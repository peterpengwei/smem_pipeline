
`define PER_H 2.5
`define PER_HH 1.25

module sim_afu_core();

	reg                             CLK_400M;
    reg                             reset_n;
    
	//---------------------------------------------------
    //reg                             spl_enable;
	reg 							core_start;
	//---------------------------------------------------
	
    reg                             spl_reset;
    
    // TX_RD request; afu_core --> afu_io
    reg                             spl_tx_rd_almostfull;
    wire                              cor_tx_rd_valid;
    wire  [57:0]                      cor_tx_rd_addr;
    wire  [5:0]                       cor_tx_rd_len;  //[licheng]useless.
    
    
    // TX_WR request; afu_core --> afu_io
    reg                             spl_tx_wr_almostfull;    
    wire                              cor_tx_wr_valid;
    wire                              cor_tx_dsr_valid;
    wire                              cor_tx_fence_valid;
    wire                              cor_tx_done_valid;
    wire  [57:0]                      cor_tx_wr_addr; 
    wire  [5:0]                       cor_tx_wr_len; 
    wire  [511:0]                     cor_tx_data;
             
    // RX_RD response; afu_io --> afu_core
    reg                             io_rx_rd_valid;
    reg [511:0]                     io_rx_data;    
                 
    // afu_csr --> afu_core; afu_id
    reg                             csr_id_valid;
    wire                              csr_id_done;    
    reg [31:0]                      csr_id_addr;
        
     // afu_csr --> afu_core; afu_ctx   
    reg                             csr_ctx_base_valid;
    reg [57:0]                      csr_ctx_base;

	reg  [63:0]	dsm_base_addr;	
	reg  [63:0] 						io_src_ptr;
	reg  [63:0] 						io_dst_ptr;
	
	initial forever #`PER_HH CLK_400M=!CLK_400M;
	
	initial begin
		CLK_400M = 1;
		reset_n = 0;
		
		//---------------------------------------------------
		//spl_enable = 0;
		core_start = 0;
		//---------------------------------------------------
		
		spl_reset = 0;
		
		spl_tx_rd_almostfull = 0;
		spl_tx_wr_almostfull = 0;    

				 
		// RX_RD response = 0; afu_io --> afu_core
		io_rx_rd_valid = 0;
		io_rx_data = 0;    
					 
		// afu_csr --> afu_core = 0; afu_id
		csr_id_valid = 0;
		csr_id_addr = 0;
			
		 // afu_csr --> afu_core = 0; afu_ctx   
		csr_ctx_base_valid = 0;
		csr_ctx_base = 0;

		dsm_base_addr = 0;	
		io_src_ptr = 0;
		io_dst_ptr = 0;
		
		
		#0.1;
			
		#`PER_H;
		#`PER_H;
		
		reset_n = 1;
		
		#`PER_H;
		#`PER_H;
		
		core_start = 1;
		
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		
		io_rx_rd_valid = 1;
		io_rx_data[480] = 1; 
		io_rx_data[457:448] = 3;
		
		#`PER_H;
		
		io_rx_rd_valid = 0;
		io_rx_data = 0;
		
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		io_rx_rd_valid = 1;
		io_rx_data = 512'h00000203030303020000020002000300010303030301030303030100000200030200020200000003010000010301010302030203020300020302010301000303;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000001020203030300030002020302000001020301030000020203020303030303010301020100;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;
		io_rx_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;
		
		io_rx_data = 512'h03020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010103030003030202020003030202020003030202020003030202020003030202020003;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;
		io_rx_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;
		
		io_rx_rd_valid = 0; #`PER_H;#`PER_H;#`PER_H;#`PER_H;
		io_rx_rd_valid = 1;
		
		io_rx_data = 512'h00000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000300;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000001000003000101000003010101000103010101000003020101000003010101000003020101;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;
		io_rx_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;
		io_rx_rd_valid = 0;
		
		#300;
		io_rx_rd_valid = 1;
		
		io_rx_data = 512'h40003001000040030040000000000000000103010400400040000000900040000000000000000000000000000000000000000000000000000000000000000000;#`PER_H;
		io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_data = 512'he8eccedcbecc0fbbe9cc8af1f5809048dfd7bb5fdefe5df6f5c3bffe3ffffe69000000002e38563c00000000265dfe18000000002e1ed23000000000362ca1fc;#`PER_H;
		io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_data = 512'h6bfa2ffe000000004ce798c5000000004ce798c5000000006bfa2ffeffc00000000000006bfa2ff9000000004ce798c5000000004ce798c5000000006bfa2ffd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h40003001000040030040000000000000000103010400400040000000900040000000000000000000000000000000000000000000000000000000000000000000;#`PER_H;
		io_rx_data = 512'h550eff5ff77db4376975d17bdfccea5988e3269e22c92f30b3f93ffcdda9fbee00000000078b380d00000000072d0e630000000006e96251000000000d90bdbf;#`PER_H;
		io_rx_data = 512'h3b373318cc38016903dff27bc00d1763339d3fa6962fefe1cfa0c0d98d6a071e000000001f51358c000000001b64c34500000000214ce72e000000002a86c281;#`PER_H;
		io_rx_data = 512'hffb3337f5637fd1df6f3807f8fdf74c7761ffb95eac16d48facfbfdc7feef435000000002507a8a3000000001fe5dfeb00000000263b379e000000002ef041d4;#`PER_H;
		io_rx_data = 512'h0412571d5c554102081c05d5c0474105c04564346113343870ecd31500afbcdf0000000010b47bd7000000001108779b0000000013d8aa3c000000001a3db452;#`PER_H;
		io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_data = 512'h1157157d740015301145110c54754154540175d537d7577205f15dfe5d5d571f000000004b29eeee000000003b3fc6850000000034b17a6100000000523969ac;#`PER_H;
		io_rx_data = 512'hdfdfdffdfd77cfeff51d7f433f7db7ff93d63e77ac963f7dd1e63f3f9b1a89bf00000000211c4ace000000001ce182ca00000000233180f3000000002c17c875;#`PER_H;
		io_rx_data = 512'hfcfda0ff4cffcf1ff4ef1c337fff0cff4c3fde4ecffdb73172b8dea48f3ffbbb0000000022b66fea000000001df0515000000000245bfefa000000002d32a74c;#`PER_H;
		io_rx_data = 512'h719779259a8bcd45cb8787fd136d81614cb5234e44f1b04f5d1577fdcbbba5cf000000004dece9a6000000003cfc0ba20000000036c1252f0000000054d3c289;#`PER_H;
		io_rx_data = 512'h555555515555555545555555555555d5555555555555555555555575cbd3e5150000000050530159000000003e3e1a9f0000000038196f4f00000000574e8c39;#`PER_H;
		
		io_rx_rd_valid = 0;
		spl_tx_rd_almostfull = 1;
		
		
		
		#150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h3202b32b08033f08cebe80b773803c3f8f7f36ee33bbb31ef90fcc8fc03ffefc0000000041736d3d000000003583de3e0000000031f437490000000049e3a33c;#`PER_H;
		io_rx_data = 512'hff0c032ac2b003f3fbc3f3fec3efeffb0ceafcac8f9fe1bc80fbefeeaeea23ea0000000041ffb8530000000035c9200500000000320661f3000000004a5254b5;#`PER_H;
		io_rx_data = 512'h67ff1dd01e748504d4655d55855835a875c75f5071ed86ca00070055c34f3b6700000000099b448d0000000008dba8e70000000009727bc500000000102e5ec7;#`PER_H;
		io_rx_data = 512'h8c7d0f4c5a864fdc73cf36f93e9d7424f416b1f715265f70df7ecddff418448d0000000009d2443f000000000912cb270000000009cc10630000000010818737;#`PER_H;
		io_rx_data = 512'h7ddcbf05e5d9d71335dc5fbfceff6fffc45bde10ffcec7bff3feff5e33ff47ad0000000060559ac100000000484410ee0000000046a31e2c0000000064798125;#`PER_H;
		io_rx_data = 512'hff67ffdd405dffff901c14731407cd1bc4e0430e3f47800a0e1d35444d43d828000000006154cecd0000000048973f600000000047072ef10000000065292562;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h03143c734765f40cda19020ff1d35fa5fc82c565f245e2c303efbad7355b9dd1000000000f78a45b000000000fbd150600000000123ae0680000000018730937;#`PER_H;
		io_rx_data = 512'h0000e90000040119040c0010ad401000d57f235c4a416d57c25954e1d15312c3000000000f91151d000000000fd12f3600000000125725ed000000001898ea40;#`PER_H;
		io_rx_data = 512'h5c100147902c801415494444d0cb0438357814ff43ed0f878006dcdc8c97b0f1000000000372bd11000000000327ca2000000000032b929500000000066844ba;#`PER_H;
		io_rx_data = 512'h7000c2c5a0d45778292507eff5db2f078463f1d04dc1234714438bae3453d5c400000000037feb9100000000033b96e400000000033cbd6c000000000689471f;#`PER_H;
		io_rx_data = 512'h00f8a033f3ceff03f0c20208ffc0cf8e8ecefff3cf0c8fbfd3033ffbfb53f0c70000000046e595820000000038e1193c0000000032fd274e000000004e620374;#`PER_H;
		io_rx_data = 512'heb2c0c0330e3f3f1b37b008bf00cfd84fcfecb6ffff06ed72bffffb3b7acbaf60000000047080fe60000000038f199b9000000003301f782000000004e7d66df;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h048fc233c288ff303ff3ecbcf43cf3b0b7e0f88fcfc0b093cfec3ff83e30c30b00000000333e4237000000002a7662ad000000002ef37a88000000003bf6be14;#`PER_H;
		io_rx_data = 512'hffeff383e98caaff48eebfcfff3bfcfffc3b032c2c81fc03383023fccc000f8b00000000334543d1000000002a7ac7d1000000002ef46f4a000000003bfe7d14;#`PER_H;
		io_rx_data = 512'hceb6014be67cfed412c4fef08202c3c1b8bdbc3cbec9fe97ff39b6a1fb537fff0000000049e7380d000000003a798f9a0000000033dfc2a10000000050fb9438;#`PER_H;
		io_rx_data = 512'h56000b33f043c07f32ef1db0fd040419766c50c0c3df27346c243fe0344c43960000000049eaf923000000003a7c475b0000000033e2ee690000000050ff1e19;#`PER_H;
		io_rx_data = 512'hf3d3ffc28ca0bcf2f2c8dcbf22803ecbbfbc6208eff2fb0e03c280aeca203fc2000000004116522900000000353a5a730000000031e5fb0c00000000498c3a58;#`PER_H;
		io_rx_data = 512'hfabe3ffcfefbe3b4ffbc7f7ced70eecbf72cc23cdf3edf31c08f0f8caf3fc5d800000000411ce5f500000000353de4610000000031e6d614000000004991c216;#`PER_H;
		
		spl_tx_rd_almostfull = 0;
		
		
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0e1393cf6c0d4e01c04c3383f514d0c0c30f3fe6dc8f2c012dacc362d7eecbc300000000253c46cf0000000020167049000000002675cdfb000000002f25256d;#`PER_H;
		io_rx_data = 512'hffff218200c3ffff70c1c785c77d4031f7444f607555dd7c0c09dce5a245555300000000253c80270000000020169ece000000002676170d000000002f2568fe;#`PER_H;
		io_rx_data = 512'h20b5630743f0f5133f0fcf7414b788fa0d54f0227f75314f6dfdb7965d97f5bd000000002668ae8900000000214462790000000027befb0b00000000306de673;#`PER_H;
		io_rx_data = 512'hd1bdcb8cf04f773d29cec18feffffd21fe3c5d3ff7afdc37fe72a667d7757c6d000000002669a464000000002144dba30000000027c009f600000000306e9403;#`PER_H;
		io_rx_data = 512'h0be3080b03df0fc3ef3d8bc2eb838be188efa80ce882702ca8ce6b8ecaabccbf000000003fc870e300000000345424550000000031a5af90000000004859de38;#`PER_H;
		io_rx_data = 512'haaec30b0fff7aaaafb837f8cea2baa3c2f23fb3effefe00dfaf23af73328fb02000000003fc9d85f000000003454f3620000000031a5e56300000000485afbdc;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h3d814ffc74bb3cc53788d1054371bbff798d35d7c6203f4f2ae8f65a70bd3c7b000000000a3e3a2e0000000009763339000000000a6aab250000000011060c74;#`PER_H;
		io_rx_data = 512'hf220f5116a81008009470ddc0d2582505c0784d333c8c89331e00dc1c91071a7000000000a3e48dc000000000976417b000000000a6ac0920000000011061e17;#`PER_H;
		io_rx_data = 512'h4557755b5557d7503f55d5d5ad00f93397cf0cffcd13958fbadb9ff7eb77cf140000000023111e19000000001e508b550000000024d3d2e3000000002d83aeaf;#`PER_H;
		io_rx_data = 512'hbffc458fdd5eff1f5b79edc35ffe47861ea3f5750cdf2b706c7732f1b075469000000000231170b0000000001e50af160000000024d437b4000000002d83e286;#`PER_H;
		io_rx_data = 512'h201941a780017055d490932055b117b4038e1101dd90e0e22f09443cf9df557f000000000f2d505e000000000f52ecf20000000011c7c227000000001811de89;#`PER_H;
		io_rx_data = 512'h642dac53dba36b95d61ba004c208bfd5b47f8052dd2c278725fc5ded83efde99000000000f2d98eb000000000f531fce0000000011c8179d0000000018122b2a;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'ha464f84210c99f73f24d23453c332c1115e28320bc0dfb5a36473ef357025c05000000001af5de22000000001814eaee000000001d246389000000002635ae67;#`PER_H;
		io_rx_data = 512'h54f1008cf7a8c3e7b1c7ffff01f11f1f51dbdc04413c1335dd900c529d08e7f0000000001af5e0c1000000001814f1fa000000001d2469b7000000002635b40e;#`PER_H;
		io_rx_data = 512'hdfaf7c7ff578740c7f19fcbec80f9a33f9fc0bde80fcd75d3e94bbc4f3fffff000000000223d2c29000000001da5c735000000002407d8c7000000002ce3365b;#`PER_H;
		io_rx_data = 512'h3fbe74e10b6e82a9f73e47cc06b12096136f3f303d0d4fcd1fdc18b83dbdb3f700000000223d471d000000001da5d7df000000002407f5b5000000002ce352cf;#`PER_H;
		io_rx_data = 512'h3b57ced710f073c974138fc3dd578ffdf24323fff34f2c3540ffdfbc6f7fd4f3000000004d73634e000000003cabe61c000000003672bb97000000005464ac7f;#`PER_H;
		io_rx_data = 512'h54b00c700d93ad401453f18f3e3ecf1f54dd874f3341455f56fe5c2f1c915502000000004d7378df000000003cabf2dd000000003672ccd2000000005464c1f2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h8b3330d5178c369d4ff3b3ea05840b4505a0505f7c505c00b7dabf0e5fcdcf4e00000000513bc351000000003eb090000000000038d3fc960000000057feef99;#`PER_H;
		io_rx_data = 512'h0cff418d898a50a447c6083cc734059ff622bc0f719e13fd1c70d9bf37cc113100000000513bc407000000003eb090730000000038d3fd370000000057fef04f;#`PER_H;
		io_rx_data = 512'h37e01403ddc121ff2869570c3135076448543e563433b7cbf3833315edf300300000000009c245a000000000090129aa0000000009b4e74500000000106adf71;#`PER_H;
		io_rx_data = 512'h769704cb8807cbdd4345f5056c00cc50ff20243c2890880c604425e13035f8040000000009c248950000000009012f7b0000000009b4ec1300000000106aee5d;#`PER_H;
		io_rx_data = 512'h3eac3efffff12ef13fd8c240f3034cc01cf3cdcf327efb42f3ff07e7133be3f4000000006023eda0000000004832028200000000468c24dc00000000645ab002;#`PER_H;
		io_rx_data = 512'h3880001cb386d2bffffbf7f33cfceacf03830f7a39e913cf7ebf97cd33bd4f1f000000006023f54600000000483205a900000000468c2a1a00000000645ab4f7;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h304cac3d5ecd1c0efeb2c7cb5b3a01ef8b1727f094803a1d01403e3e52aaab870000000012fe9bc200000000125cdc34000000001584b701000000001d1ec089;#`PER_H;
		io_rx_data = 512'hac9217933d56c4d8504715d35d4f1c80ddc940a1d6e58801915b8144413b5c720000000012fe9be600000000125cdc52000000001584b717000000001d1ec0b1;#`PER_H;
		io_rx_data = 512'hf7ffd55c3ff7ffff551f3cfd0f470f31f3943f5afdf430b401d7443d15908f9e00000000037bee2a0000000003376f3200000000033805f600000000067f7c2e;#`PER_H;
		io_rx_data = 512'h51f14f25fff0d41433ffffff03b43bc4a90ffd80eb58113a1f7210a627c1c7c000000000037bf723000000000337704100000000033807be00000000067f7f5e;#`PER_H;
		io_rx_data = 512'hcf7eebfa22002bcbc3f33eac22083f0c2822eaa72b9c2eba30e835e9ab82aaba0000000046de25ff0000000038dd43db0000000032fbdb86000000004e5c85a0;#`PER_H;
		io_rx_data = 512'hb10f332f2bcc73f7ca80f2003cfbef7a3fcf0ff3886ef8c3e3ef28f882bcb0ca0000000046de27100000000038dd44cd0000000032fbdba1000000004e5c8682;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'habbe5d0471f9aaa87bb3d03b7d7de581b26542aea958000dcb6332d888500140000000001de284e3000000001a6c592d0000000020082ed5000000002927da1b;#`PER_H;
		io_rx_data = 512'habbe5d0471f9aaa87bb3d03b7d7de581b26542aea958000dcb6332d888500140000000001de284e3000000001a6c592d0000000020082ed5000000002927da1b;#`PER_H;
		io_rx_data = 512'h559c301255555154555555555d65d794addb555d53f4d94d374373a687c9561d0000000049e9c2b0000000003a7b907f0000000033e1f2860000000050fe09cb;#`PER_H;
		io_rx_data = 512'h5555573515455555d4e568f5f55695ff5e15855d95195774597567295555d5d50000000049e9c34d000000003a7b90d10000000033e1fa340000000050fe0a2e;#`PER_H;
		io_rx_data = 512'h3e2bbb230ae0a8be303b0a0e0ae1bf3c1680aaaaaa28a2aaaaebaaaa3aa8bfaa000000004115087500000000353972780000000031e5c35300000000498ace40;#`PER_H;
		io_rx_data = 512'h08fe080b08b822e8aaca0bbdeea90a2eb080a83082cbe380a08ab08ebe2cbabe00000000411508af00000000353972ee0000000031e5c35900000000498ace8a;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5881d1110870100cb33d9030fcb2cf4102a0e03f001334c015d05e1c000003e20000000008f235c400000000084d9fb8000000000892851b000000000f557f69;#`PER_H;
		io_rx_data = 512'h5881d1110870100cb33d9030fcb2cf4102a0e03f001334c015d05e1c000003e20000000008f235c400000000084d9fb8000000000892851b000000000f557f69;#`PER_H;
		io_rx_data = 512'hb0555ce775e55554d5975d7f555d141e55555555755955558f55a4715515d7e30000000026695920000000002144b7810000000027bfb2c300000000306e5f1c;#`PER_H;
		io_rx_data = 512'h700015555d5574553555d0755d5759555555515555554b5555555555575d55550000000026695982000000002144b7b60000000027bfb96f00000000306e5f59;#`PER_H;
		io_rx_data = 512'h3cc2f0f2000c083032000c43b8003cc00020a008a0f02003000e2000c0c2b000000000003fc82243000000003453e7b90000000031a5a18e0000000048598f76;#`PER_H;
		io_rx_data = 512'h35a30c8c013b383fa2c0b8b220b880a8d8802ffb2bc822cb2cc0fc00fe02cc3a000000003fc8225a000000003453e7ca0000000031a5a18f0000000048598fcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h4cc6461d52984f87c0a44d9db4770809275097512342adc3fbaaa8b0aaaaaab9000000001a761c3c0000000017be2b39000000001c9061750000000025c80c16;#`PER_H;
		io_rx_data = 512'h4cc6461d52984f87c0a44d9db4770809275097512342adc3fbaaa8b0aaaaaab9000000001a761c3c0000000017be2b39000000001c9061750000000025c80c16;#`PER_H;
		io_rx_data = 512'h555155755555555517515575525573d555b1560cd55d9955bf77c55545d55357000000002311584e000000001e50a4b40000000024d417f0000000002d83cd8e;#`PER_H;
		io_rx_data = 512'h5f55649dda4e55e554ad9b415570551555d5565654d55555557173555550555500000000231158ad000000001e50a4db0000000024d41e2a000000002d83cdce;#`PER_H;
		io_rx_data = 512'h154cdeecfe3fbffdb8fffdfefbf5ff9dffffef35f7cfffffffffcff5fff0fbff000000000f2d4165000000000f52d7fc0000000011c7ad9a000000001811c885;#`PER_H;
		io_rx_data = 512'h154cdeecfe3fbffdb8fffdfefbf5ff9dffffef35f7cfffffffffcff5fff0fbff000000000f2d4165000000000f52d7fc0000000011c7ad9a000000001811c885;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hc13c3528786c40034075322d449945524ef2f5200d56f9051c5a0f120142512d0000000008251c370000000007a19c8300000000079b297f000000000e6629c7;#`PER_H;
		io_rx_data = 512'hc13c3528786c40034075322d449945524ef2f5200d56f9051c5a0f120142512d0000000008251c370000000007a19c8300000000079b297f000000000e6629c7;#`PER_H;
		io_rx_data = 512'h10013c03800001010008000005020000000000000a000000255000351003d00000000000223d409c000000001da5d37c000000002407eda4000000002ce34644;#`PER_H;
		io_rx_data = 512'h055401348000020304000000001550001501450c15502011000030c50000000200000000223d40c3000000001da5d39a000000002407ee24000000002ce34b7f;#`PER_H;
		io_rx_data = 512'hdff73ef0ffffcfd4fff7cff27ffff7fffffefff0ffc7effffffc3ffffeebffff000000004d735d6f000000003cabe391000000003672b8f4000000005464a90c;#`PER_H;
		io_rx_data = 512'hdff73ef0ffffcfd4fff7cff27ffff7fffffefff0ffc7effffffc3ffffeebffff000000004d735d6f000000003cabe391000000003672b8f4000000005464a90c;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'hb00000000000000000014c0c43f0023008078fcc1070000400150000459000000000000009c2478f0000000009012e5f0000000009b4ea8500000000106ae58d;#`PER_H;
		io_rx_data = 512'h0044f0002400010cc000805000caa00a1321008903aa000000007000000000000000000009c247c50000000009012e780000000009b4eaae00000000106aea95;#`PER_H;
		io_rx_data = 512'h822a2baa062aaa8ab8b21ab8b09eb9aaead6aebeaaeaa2abab8a6ae8aaaaae7a000000006023ebb4000000004832007d00000000468c23f000000000645aaedf;#`PER_H;
		io_rx_data = 512'h822a2baa062aaa8ab8b21ab8b09eb9aaead6aebeaaeaa2abab8a6ae8aaaaae7a000000006023ebb4000000004832007d00000000468c23f000000000645aaedf;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'h0003e03f5ffffffcc7033efffff3eefff0ffd3ffff7ffff0000fbf0ffcce03d200000000037bf05d0000000003376fd200000000033806fc00000000067f7e55;#`PER_H;
		io_rx_data = 512'hfff5ffffcf7fff9ff3df8fffffb73fffffff07ff7fffffffffdfeffffff3ffff00000000037bf4d80000000003376fe8000000000338072e00000000067f7e92;#`PER_H;
		io_rx_data = 512'haaaa62abaaaaaaa8aaa82aaa0095aa8aa82aa2aaaaa8aaeaaaaaaaaaaaaaaaaa0000000046de25c10000000038dd427d0000000032fbdb71000000004e5c8551;#`PER_H;
		io_rx_data = 512'haaaa62abaaaaaaa8aaa82aaa0095aa8aa82aa2aaaaa8aaeaaaaaaaaaaaaaaaaa0000000046de25c10000000038dd427d0000000032fbdb71000000004e5c8551;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'he839335eaf56bf785c75d47ac7ddace52efdf3dd4ca45271388104c7702da1b3000000005fb7194c0000000047fcfe3a000000004648c2230000000063fed5d7;#`PER_H;
		io_rx_data = 512'h55555d555555555557d555555555d5555555555555571655555555555555555d0000000049e9c300000000003a7b90ac0000000033e1f44b0000000050fe0a09;#`PER_H;
		io_rx_data = 512'h5555555f545455555d55a9545755557d5d5555d5555595555555715555d555f50000000049e9c31f000000003a7b90b40000000033e1f8960000000050fe0a17;#`PER_H;
		io_rx_data = 512'haaaaaa8aaa6aaea8aaaaaaaaaaaaaaaa4aaaaaaa9aaa8aaaab8aaaaaaaaaaaaa000000004115086500000000353971aa0000000031e5c34f00000000498ace22;#`PER_H;
		io_rx_data = 512'haaaaaa8aaa6aaea8aaaaaaaaaaaaaaaa4aaaaaaa9aaa8aaaab8aaaaaaaaaaaaa000000004115086500000000353971aa0000000031e5c34f00000000498ace22;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h34c0f03fbd1044485f00594155df3c48099fd1fbff1f0cbf4acfed0c7973933b000000005fb719200000000047fcfe2c000000004648c2050000000063fed5af;#`PER_H;
		io_rx_data = 512'he839335eaf56bf785c75d47ac7ddace52efdf3dd4ca45271388104c7702da1b3000000005fb7194c0000000047fcfe3a000000004648c2230000000063fed5d7;#`PER_H;
		io_rx_data = 512'h25155555555555d1555555555555555b455da5555555555575551555545555570000000026695942000000002144b7950000000027bfb3f900000000306e5f30;#`PER_H;
		io_rx_data = 512'h55555575545595545005455775c41ffd7555555555555c75555579d5555555550000000026695952000000002144b7a60000000027bfb84600000000306e5f42;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h3c855c87f43c93b307e77ef4b1470c20a6aa9aa7b722aaaaba5379d8fbc3c511000000005fb718fe0000000047fcfe07000000004648c1ea0000000063fed591;#`PER_H;
		io_rx_data = 512'he839335eaf56bf785c75d47ac7ddace52efdf3dd4ca45271388104c7702da1b3000000005fb7194c0000000047fcfe3a000000004648c2230000000063fed5d7;#`PER_H;
		io_rx_data = 512'h55a955551555555555555054d56a7455555a5d45555555555555155555555555000000002311586e000000001e50a4c20000000024d41925000000002d83cdab;#`PER_H;
		io_rx_data = 512'h9d5555555555575553554555557d55555555e5555555555555515c55555555e70000000023115885000000001e50a4cf0000000024d41cef000000002d83cdbd;#`PER_H;
		io_rx_data = 512'hdcf9507fffffcf3ffffffffffffffdffeffcffffffefffffffffff3ffdffffcf000000000f2d40f7000000000f52d7f90000000011c7ad93000000001811c87d;#`PER_H;
		io_rx_data = 512'hdcf9507fffffcf3ffffffffffffffdffeffcffffffefffffffffff3ffdffffcf000000000f2d40f7000000000f52d7f90000000011c7ad93000000001811c87d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hc606d976a0cd0767f63374f35d1fe3719ecf07fdcd2e0733f761507fc9324ce8000000005fb718680000000047fcfdca000000004648c18e0000000063fed540;#`PER_H;
		io_rx_data = 512'he839335eaf56bf785c75d47ac7ddace52efdf3dd4ca45271388104c7702da1b3000000005fb7194c0000000047fcfe3a000000004648c2230000000063fed5d7;#`PER_H;
		io_rx_data = 512'h000800001000044000007010000008000000040054000014450dce040008104000000000223d40a7000000001da5d385000000002407edcc000000002ce34708;#`PER_H;
		io_rx_data = 512'h0c030010000008000000400000010004000001500480c001001000000000051000000000223d40b4000000001da5d390000000002407ee05000000002ce34ab7;#`PER_H;
		io_rx_data = 512'hffffffffffcfffeffffffffff7ffffdfffeefffffffffffffffcfffffffff7ff000000004d735cf7000000003cabe38e000000003672b8f1000000005464a90a;#`PER_H;
		io_rx_data = 512'hffffffffffcfffeffffffffff7ffffdfffeefffffffffffffffcfffffffff7ff000000004d735cf7000000003cabe38e000000003672b8f1000000005464a90a;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hc606d976a0cd0767f63374f35d1fe3719ecf07fdcd2e0733f761507fc9324ce8000000005fb718680000000047fcfdca000000004648c18e0000000063fed540;#`PER_H;
		io_rx_data = 512'hcdef55fb78bf32b3000c82fc3ceb8000fcdf0df6fb48fa7f593c72e8d9c10fe7000000005fb71f7f0000000047fd04f3000000004648c4190000000063fed975;#`PER_H;
		io_rx_data = 512'h010000300060000000000c0008000000000000000000000000000000c00c00000000000009c247a20000000009012e6f0000000009b4ea9600000000106ae659;#`PER_H;
		io_rx_data = 512'h00000001000000080300001000000000010000003c3000003000000000c00c030000000009c247bc0000000009012e720000000009b4eaa000000000106ae9b2;#`PER_H;
		io_rx_data = 512'haaaaaaaaa2aaaabaaa0faa8aaaa96aaaaaaaabaaaa9a2eaaab83caaa8bb2abaa000000006023eba9000000004832001500000000468c23ed00000000645aaed5;#`PER_H;
		io_rx_data = 512'haaaaaaaaa2aaaabaaa0faa8aaaa96aaaaaaaabaaaa9a2eaaab83caaa8bb2abaa000000006023eba9000000004832001500000000468c23ed00000000645aaed5;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hebeefecd2f7d8c45ae06eb124bc8ffd425f6945d5cc4ff3ffea7d037d9b320ff000000005fb70f130000000047fcf3d2000000004648bd850000000063fecf96;#`PER_H;
		io_rx_data = 512'h4f318ff5b73cd3f0e439436bfcfedb2bf3de00242633c373469feffcfb830e37000000005fb726c40000000047fd071f000000004648c94e0000000063fedccf;#`PER_H;
		io_rx_data = 512'hfffff1ffefffffffffffff53dfdffffff7ff77fffff7ffffdffc3fffffffffff00000000037bf11a0000000003376fe0000000000338070b00000000067f7e7b;#`PER_H;
		io_rx_data = 512'hfffffffdfdffffffcffffff7bff70fffffffdfc3fff7ffff3fdbff55ffcfffff00000000037bf46c0000000003376fe6000000000338072300000000067f7e8b;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hd792403c83f0d5f400fdbccfffffcd20397f550b3ddd1ddd2d35e780d7bf03f7000000005fb6dd060000000047fcc3ca00000000464893240000000063feab0c;#`PER_H;
		io_rx_data = 512'h4f318ff5b73cd3f0e439436bfcfedb2bf3de00242633c373469feffcfb830e37000000005fb726c40000000047fd071f000000004648c94e0000000063fedccf;#`PER_H;
		io_rx_data = 512'h5555555555f555555555555555555d595554d555555555415f5555555d5555550000000049e9c306000000003a7b90ad0000000033e1f4c30000000050fe0a0a;#`PER_H;
		io_rx_data = 512'h5577555555545555559557555d55555551941555d95555d651555551555555550000000049e9c319000000003a7b90b00000000033e1f8260000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa2aa2aa8aaaaaaaaaaaaaaaaaaa0000000041150865000000003539712d0000000031e5c34f00000000498ace1f;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa2aa2aa8aaaaaaaaaaaaaaaaaaa0000000041150865000000003539712d0000000031e5c34f00000000498ace1f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hff68489fdbf0c925040d0b3fbf97ca0f6f2ece0d38ce5a1cfffcbf0d2386011f000000005fb2c81e0000000047faf410000000004645fd6f0000000063fbbee3;#`PER_H;
		io_rx_data = 512'hbff7fafd396f183f7133dd7ba77fd0ab6eba254347e54112beff54674cf77f7d000000005fba0a690000000047fe21e400000000464abaaf000000006400ab84;#`PER_H;
		io_rx_data = 512'h5595555545555555155565555555555555555555555555555555555555555555000000002669594b000000002144b79e0000000027bfb4e000000000306e5f37;#`PER_H;
		io_rx_data = 512'h55515755555555555755555555575d5655555195555595555555555575555555000000002669594d000000002144b7a30000000027bfb7d000000000306e5f40;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfdfcfffefffcfffdbfec43f6bff5f2b1c6fb73dfff3fbfbecffc33ffdefe9e0d000000005faa0dc80000000047f7094000000000464112920000000063f4de66;#`PER_H;
		io_rx_data = 512'h73d3ccdd2b73ec9c7743cfefbb37bfddd3f4f1ef331755c6cc7bc77f92fd40d8000000005fd294c90000000048092cef000000004657a06f00000000641256d9;#`PER_H;
		io_rx_data = 512'h5555555555555555c55515b555555745665555d55fd55555555555555d5515550000000023115871000000001e50a4ca0000000024d41993000000002d83cdb2;#`PER_H;
		io_rx_data = 512'h55d155555515d555555555555d5555555555555555555557555d5655555555550000000023115880000000001e50a4ce0000000024d41c77000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h4bff5c3fbff71f2d7b13f3f06f037ff2d3c3b7fecff3c9f44cf7fe278fc754fc000000005f5f923c0000000047d2edba000000004614d9dc0000000063abf6ae;#`PER_H;
		io_rx_data = 512'h73d3ccdd2b73ec9c7743cfefbb37bfddd3f4f1ef331755c6cc7bc77f92fd40d8000000005fd294c90000000048092cef000000004657a06f00000000641256d9;#`PER_H;
		io_rx_data = 512'h4000000119400030300054000014c1000000000030000600000101000010300000000000223d40ab000000001da5d389000000002407edde000000002ce3476e;#`PER_H;
		io_rx_data = 512'h0000100010040000003800000001010000400a0300c10100000000000010000000000000223d40b1000000001da5d38d000000002407edfc000000002ce34a46;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h01d565d96bc4fb55bcdf26551f5f7d51f7bde5d714ba55ea6167526d9fd77d52000000005e69721f00000000477bf8560000000045a642810000000063057d8a;#`PER_H;
		io_rx_data = 512'hff67ffdd405dffff901c14731407cd1bc4e0430e3f47800a0e1d35444d43d828000000006154cecd0000000048973f600000000047072ef10000000065292562;#`PER_H;
		io_rx_data = 512'h000000000000000000004c0000000003000000000302000c0000000f00030c000000000009c247a60000000009012e710000000009b4ea9800000000106ae6d1;#`PER_H;
		io_rx_data = 512'h00000001000000080300001000000000010000003c3000003000000000c00c030000000009c247bc0000000009012e720000000009b4eaa000000000106ae9b2;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h01d565d96bc4fb55bcdf26551f5f7d51f7bde5d714ba55ea6167526d9fd77d52000000005e69721f00000000477bf8560000000045a642810000000063057d8a;#`PER_H;
		io_rx_data = 512'h6bfa2ffe000000004ce798c5000000004ce798c5000000006bfa2ffeffc00000000000006bfa2ff9000000004ce798c5000000004ce798c5000000006bfa2ffd;#`PER_H;
		io_rx_data = 512'hfffffffdffffff3ff3ffffffffd7ffffffcffffff7ffffffffffffffffffdfef00000000037bf18b0000000003376fe1000000000338071500000000067f7e7f;#`PER_H;
		io_rx_data = 512'hfffffffff7cbfffffffffffffffffffffffffffffffff3cffffffbdcffffffff00000000037bf3f40000000003376fe4000000000338072100000000067f7e87;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_data = 512'h6bfa2ffe000000004ce798c5000000004ce798c5000000006bfa2ffeffc00000000000006bfa2ff9000000004ce798c5000000004ce798c5000000006bfa2ffd;#`PER_H;
		io_rx_data = 512'h55515555555555555555555595555554515555555555555555d55555b55555550000000049e9c30d000000003a7b90ae0000000033e1f5380000000050fe0a0d;#`PER_H;
		io_rx_data = 512'h5555555555555555755555dd5555555555555555555557555555d5555555d5550000000049e9c313000000003a7b90b00000000033e1f7ac0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5595555545555555155565555555555555555555555555555555555555555555000000002669594b000000002144b79e0000000027bfb4e000000000306e5f37;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555515555555d577555555555551555755555555555f55195550000000023115879000000001e50a4cd0000000024d41a04000000002d83cdb6;#`PER_H;
		io_rx_data = 512'h55d155555515d555555555555d5555555555555555555557555d5655555555550000000023115880000000001e50a4ce0000000024d41c77000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0100000000000000200040004400c0004400000000000000040004000001000000000000223d40b0000000001da5d38b000000002407eded000000002ce347d8;#`PER_H;
		io_rx_data = 512'h0000100010040000003800000001010000400a0300c10100000000000010000000000000223d40b1000000001da5d38d000000002407edfc000000002ce34a46;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffdffffff3ff3ffffffffd7ffffffcffffff7ffffffffffffffffffdfef00000000037bf18b0000000003376fe1000000000338071500000000067f7e7f;#`PER_H;
		io_rx_data = 512'hfffffffff7cbfffffffffffffffffffffffffffffffff3cffffffbdcffffffff00000000037bf3f40000000003376fe4000000000338072100000000067f7e87;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_data = 512'haea2aaaaaa8aaaaaaaaabaaaabaaaaaaaaaaaaaaaaaaaaaeaaaaabaaaaaaaaea0000000046de25bb0000000038dd42050000000032fbdb71000000004e5c854f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h55515555555555555555555595555554515555555555555555d55555b55555550000000049e9c30d000000003a7b90ae0000000033e1f5380000000050fe0a0d;#`PER_H;
		io_rx_data = 512'h5555555555555555755555dd5555555555555555555557555555d5555555d5550000000049e9c313000000003a7b90b00000000033e1f7ac0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555515555555d577555555555551555755555555555f55195550000000023115879000000001e50a4cd0000000024d41a04000000002d83cdb6;#`PER_H;
		io_rx_data = 512'h55d155555515d555555555555d5555555555555555555557555d5655555555550000000023115880000000001e50a4ce0000000024d41c77000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hfffff7dffffffffffcfffd007fffffffffffffffffffffffffffffffffffffff000000000f2d4080000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0100000000000000200040004400c0004400000000000000040004000001000000000000223d40b0000000001da5d38b000000002407eded000000002ce347d8;#`PER_H;
		io_rx_data = 512'h0000100010040000003800000001010000400a0300c10100000000000010000000000000223d40b1000000001da5d38d000000002407edfc000000002ce34a46;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hffffcfffffffffffffffffffffff7ffffffffffffcffffffeffbffffffffffff000000004d735c7c000000003cabe38c000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffdffffff3ff3ffffffffd7ffffffcffffff7ffffffffffffffffffdfef00000000037bf18b0000000003376fe1000000000338071500000000067f7e7f;#`PER_H;
		io_rx_data = 512'hfffffffff7cbfffffffffffffffffffffffffffffffff3cffffffbdcffffffff00000000037bf3f40000000003376fe4000000000338072100000000067f7e87;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h55515555555555555555555595555554515555555555555555d55555b55555550000000049e9c30d000000003a7b90ae0000000033e1f5380000000050fe0a0d;#`PER_H;
		io_rx_data = 512'h5555555555555555755555dd5555555555555555555557555555d5555555d5550000000049e9c313000000003a7b90b00000000033e1f7ac0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55d155555515d555555555555d5555555555555555555557555d5655555555550000000023115880000000001e50a4ce0000000024d41c77000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0100000000000000200040004400c0004400000000000000040004000001000000000000223d40b0000000001da5d38b000000002407eded000000002ce347d8;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaa8aaaaaaeaa9eaaaaaa8aaaaaaaeaeaaaabaaaae9a2aaaaeaaaaaaaaaaaba000000006023eba1000000004831ffa200000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555595555055555555555555555555555555555555555555555515555000000002669594d000000002144b7a20000000027bfb75400000000306e5f3d;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff000000000f2d4000000000000f52d7f90000000011c7ad8f000000001811c878;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffffbfeffffffffffffffffffffffffffffffffff000000004d735bfe000000003cabe38a000000003672b8f0000000005464a908;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0040000000c0000000000000300000000000f0000c00000100000000000000300000000009c247ae0000000009012e720000000009b4ea9900000000106ae747;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000006023eba0000000004831ff2300000000468c23eb00000000645aaed2;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_data = 512'haaaaaaaaaaaaaaaaaaaaaaaaaaa8aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000000046de25bb0000000038dd41860000000032fbdb71000000004e5c854e;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_data = 512'haaaaaabaaaaa2a2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000000004115086400000000353970b00000000031e5c34f00000000498ace1d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555555555595555555555d55555555555555555555555555555555555000000002669594c000000002144b7a10000000027bfb6d600000000306e5f3d;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010003000000000009c247b40000000009012e720000000009b4ea9b00000000106ae7bf;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555555555595555555555d55555555555555555555555555555555555000000002669594c000000002144b7a10000000027bfb6d600000000306e5f3d;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010003000000000009c247b40000000009012e720000000009b4ea9b00000000106ae7bf;#`PER_H;
		io_rx_data = 512'h0000000c00000010010000000000000003c03c01000000c300000000000000000000000009c247b50000000009012e720000000009b4ea9d00000000106ae93c;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5455555555555555555555555555555555555555555555555555555555515595000000002669594b000000002144b7a00000000027bfb55c00000000306e5f39;#`PER_H;
		io_rx_data = 512'h5555555555555555595555555555d55555555555555555555555555555555555000000002669594c000000002144b7a10000000027bfb6d600000000306e5f3d;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'h545611b05eb43a550ffdc3c0fc5556a89d2a0c55fcd5d44681e1a3704d33cfc0000000001100799e000000001134e87100000000140d342a000000001abb7347;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010003000000000009c247b40000000009012e720000000009b4ea9b00000000106ae7bf;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000400000000000000000000009c247b50000000009012e720000000009b4ea9c00000000106ae8bd;#`PER_H;
		io_rx_data = 512'h545611b05eb43a550ffdc3c0fc5556a89d2a0c55fcd5d44681e1a3704d33cfc0000000001100799e000000001134e87100000000140d342a000000001abb7347;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'h0109b13fc324d04ff0303f21af54919c0ef141034018320dd0b113d0a5e1700f000000001100793d000000001134e84100000000140d33cd000000001abb72b5;#`PER_H;
		io_rx_data = 512'h3afc5c042461030531a12106b247c21041c1cec527389c802d9e9c24c81507000000000011007a19000000001134e8c100000000140d34be000000001abb73e8;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'h5d29483fc762bc501cd43cf0f1377810a231050bf23385dac08b074c17c0d6100000000011007755000000001134e73600000000140d3252000000001abb6fa3;#`PER_H;
		io_rx_data = 512'h0c09f300f003c8303347a307d1e00e0033601c609911cf7fd4595dc30f36b1dc0000000011007c19000000001134ea1900000000140d384c000000001abb7702;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555555555555555555555555575555555000000002669594b000000002144b7a10000000027bfb5d900000000306e5f3b;#`PER_H;
		io_rx_data = 512'h5555555555555555595555555555d55555555555555555555555555555555555000000002669594c000000002144b7a10000000027bfb6d600000000306e5f3d;#`PER_H;
		io_rx_data = 512'h5d29483fc762bc501cd43cf0f1377810a231050bf23385dac08b074c17c0d6100000000011007755000000001134e73600000000140d3252000000001abb6fa3;#`PER_H;
		io_rx_data = 512'h50240688ec03d9a84766522c4820476102b0b111ce20cdc5c200c3ee593fcf33000000001100865b000000001134ef8300000000140d44c5000000001abb8e5d;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'h5d29483fc762bc501cd43cf0f1377810a231050bf23385dac08b074c17c0d6100000000011007755000000001134e73600000000140d3252000000001abb6fa3;#`PER_H;
		io_rx_data = 512'h705e101d300733d58085109f82c44f1083446e3793b50a2fe179f7f23ef03cf3000000001100b92200000000113513f300000000140d78c2000000001abbd829;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'h8cc0e421045f6f1000c201cfbe8073c48f61ced193443f2f13555a430c4f55440000000010ffd2bb0000000011347fae00000000140caf40000000001aba9257;#`PER_H;
		io_rx_data = 512'h705e101d300733d58085109f82c44f1083446e3793b50a2fe179f7f23ef03cf3000000001100b92200000000113513f300000000140d78c2000000001abbd829;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010003000000000009c247b40000000009012e720000000009b4ea9b00000000106ae7bf;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000400000000000000000000009c247b50000000009012e720000000009b4ea9c00000000106ae8bd;#`PER_H;
		io_rx_data = 512'h00c013019221049642685990811423c54744a466087122014511b7dd8c20f80e0000000010fe4198000000001133743900000000140b6212000000001ab7e81d;#`PER_H;
		io_rx_data = 512'hb8801c38054440b0dd08300d7bfa917f15d1f17e53ad6b10010cc18015c7d2f50000000011026aad000000001136365600000000140ee588000000001abdf9f5;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_data = 512'h1403e3075cf170d51140488760d34b9d00e10b00100c003102c54010c0d92c780000000010f5966600000000112dd5dc000000001404b2bd000000001aaa6701;#`PER_H;
		io_rx_data = 512'h12222f31f044e043008248c310829e81e73cc409a1c4c1084378c03cb4783a0e00000000110a7b6100000000113be0fe0000000014154049000000001aca17d8;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_data = 512'h0412571d5c554102081c05d5c0474105c04564346113343870ecd31500afbcdf0000000010b47bd7000000001108779b0000000013d8aa3c000000001a3db452;#`PER_H;
		io_rx_data = 512'h00000310000002cc0c0010004804303020030000ec8e8fed03a3049a92c38a23000000001154daa70000000011690491000000001448d06d000000001b32b9db;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555555555555555555555555575555555000000002669594b000000002144b7a10000000027bfb5d900000000306e5f3b;#`PER_H;
		io_rx_data = 512'h5555555555555555595555555555d55555555555555555555555555555555555000000002669594c000000002144b7a10000000027bfb6d600000000306e5f3d;#`PER_H;
		io_rx_data = 512'h0412571d5c554102081c05d5c0474105c04564346113343870ecd31500afbcdf0000000010b47bd7000000001108779b0000000013d8aa3c000000001a3db452;#`PER_H;
		io_rx_data = 512'h75dfdddd77d7fdfffdd5d1d5cf7d75d33fffd11ffffcddfffff0fffcffffffff0000000012d5eb6d000000001239b3d4000000001558edbc000000001ce5ff03;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555555555555555555555555555555515555555555555555555515555555000000002311587f000000001e50a4ce0000000024d41a7a000000002d83cdb9;#`PER_H;
		io_rx_data = 512'h55555555555555555555555555555555555555555555555555555555555555550000000023115880000000001e50a4ce0000000024d41bf7000000002d83cdbb;#`PER_H;
		io_rx_data = 512'h0412571d5c554102081c05d5c0474105c04564346113343870ecd31500afbcdf0000000010b47bd7000000001108779b0000000013d8aa3c000000001a3db452;#`PER_H;
		io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000000000000000000000000000000000000000000000000000000000000041000000000223d40b1000000001da5d38c000000002407edf6000000002ce3484d;#`PER_H;
		io_rx_data = 512'h000020000000000000000001000000044000000000000000000000000000004000000000223d40b1000000001da5d38c000000002407edf8000000002ce349cb;#`PER_H;
		io_rx_data = 512'h40003001000040030040000000000000000103010400400040000000900040000000000000000000000000000000000000000000000000000000000000000000;#`PER_H;
		io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000010003000000000009c247b40000000009012e720000000009b4ea9b00000000106ae7bf;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000400000000000000000000009c247b50000000009012e720000000009b4ea9c00000000106ae8bd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfffffffffffffffffdff7ffff4ffffffffffffffdff7ffcfffffdfffffb7ffcf00000000037bf2020000000003376fe2000000000338071a00000000067f7e82;#`PER_H;
		io_rx_data = 512'hfffffffffffffffffffffffffff3fffeffffffffffffffffffffffffffffffff00000000037bf3760000000003376fe3000000000338072100000000067f7e86;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h5555555551555555555555555755555555555d555555555555575555555555550000000049e9c30f000000003a7b90b00000000033e1f5b10000000050fe0a10;#`PER_H;
		io_rx_data = 512'h55555555d55555555555555555555555555555555555555555555555555555550000000049e9c312000000003a7b90b00000000033e1f72d0000000050fe0a11;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_data = 512'h61457025043027c0040fccdd94cd999815dfdbcd7c7489bd275557736530517000000000110079be000000001134e88400000000140d3453000000001abb736b;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000000000000000000000000000000000000000000000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598ccd;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h001000a000080000003000000000000000000000002000000000000000000000000000003fc82222000000003453e7860000000031a5a18b0000000048598dcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000000a00002c000000000080000080a000000008000008000282000000c00000000003fc82220000000003453e77a0000000031a5a18b0000000048598c5b;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h002000000000808000000202000000000040210000203000020e000000000200000000003fc82223000000003453e78a0000000031a5a18c0000000048598e47;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h000020000200b30080a802002000020302000000800000080080202023000002000000003fc8221c000000003453e7680000000031a5a18b0000000048598bf1;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000280a0003800830000020000c0c8a800080002000c280000020c00800080000000003fc82216000000003453e7560000000031a5a18b0000000048598b89;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000280a0003800830000020000c0c8a800080002000c280000020c00800080000000003fc82216000000003453e7560000000031a5a18b0000000048598b89;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000280a0003800830000020000c0c8a800080002000c280000020c00800080000000003fc82216000000003453e7560000000031a5a18b0000000048598b89;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000280a0003800830000020000c0c8a800080002000c280000020c00800080000000003fc82216000000003453e7560000000031a5a18b0000000048598b89;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00000280a0003800830000020000c0c8a800080002000c280000020c00800080000000003fc82216000000003453e7560000000031a5a18b0000000048598b89;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00280000a2a00820800000000000002a00c0800a000028300ac82030a0200000000000003fc82212000000003453e73d0000000031a5a18b0000000048598b26;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00280000a2a00820800000000000002a00c0800a000028300ac82030a0200000000000003fc82212000000003453e73d0000000031a5a18b0000000048598b26;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00280000a2a00820800000000000002a00c0800a000028300ac82030a0200000000000003fc82212000000003453e73d0000000031a5a18b0000000048598b26;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00820000020000000c033000a02a802a0000330808802000802e202042282008000000003fc8220c000000003453e7230000000031a5a18a0000000048598ac7;#`PER_H;
		io_rx_data = 512'h000000038f000003cc00000a0020000cc3a80000008002000000000820000080000000003fc82225000000003453e7940000000031a5a18e0000000048598eb9;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00820000020000000c033000a02a802a0000330808802000802e202042282008000000003fc8220c000000003453e7230000000031a5a18a0000000048598ac7;#`PER_H;
		io_rx_data = 512'h202a0c328abff0008000ffff000000000f3022000002080000080228f8a808e8000000003fc8222e000000003453e7a00000000031a5a18e0000000048598f24;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h00820000020000000c033000a02a802a0000330808802000802e202042282008000000003fc8220c000000003453e7230000000031a5a18a0000000048598ac7;#`PER_H;
		io_rx_data = 512'h202a0c328abff0008000ffff000000000f3022000002080000080228f8a808e8000000003fc8222e000000003453e7a00000000031a5a18e0000000048598f24;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0080808268c3c200280002488000000220200002a800a000000c0002a2800000000000003fc82204000000003453e6ec0000000031a5a1860000000048598a0a;#`PER_H;
		io_rx_data = 512'h202a0c328abff0008000ffff000000000f3022000002080000080228f8a808e8000000003fc8222e000000003453e7a00000000031a5a18e0000000048598f24;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h0000400a00000000004202a8c00000c3000b28b00c0c82b8c0300e0806800c2c000000003fc821f7000000003453e6d80000000031a5a18300000000485989ae;#`PER_H;
		io_rx_data = 512'h3cc2f0f2000c083032000c43b8003cc00020a008a0f02003000e2000c0c2b000000000003fc82243000000003453e7b90000000031a5a18e0000000048598f76;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hae000000000c000333020300c008000c202efcc0cbb03288122000020cafc008000000003fc821e2000000003453e6c50000000031a5a1820000000048598957;#`PER_H;
		io_rx_data = 512'h3cc2f0f2000c083032000c43b8003cc00020a008a0f02003000e2000c0c2b000000000003fc82243000000003453e7b90000000031a5a18e0000000048598f76;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hcc880888c03ea080ce808c833efcb282deaa246c0a8aab0f00ec338effb82000000000003fc821b1000000003453e67f0000000031a5a17e00000000485988d2;#`PER_H;
		io_rx_data = 512'h35a30c8c013b383fa2c0b8b220b880a8d8802ffb2bc822cb2cc0fc00fe02cc3a000000003fc8225a000000003453e7ca0000000031a5a18f0000000048598fcd;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hcc880888c03ea080ce808c833efcb282deaa246c0a8aab0f00ec338effb82000000000003fc821b1000000003453e67f0000000031a5a17e00000000485988d2;#`PER_H;
		io_rx_data = 512'hbfea23fffcafe3cf26e0eff20db3bacaccf8ebcb2a8e92f0fea2b00200b028be000000003fc823a3000000003453e9ee0000000031a5a1bd0000000048599232;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hbdef80fb33fff00cfa2332ae30eefcfc208688333aafc0e3e8ab0238aaaa8e30000000003fc81bbc000000003453e3560000000031a5a11c00000000485984d2;#`PER_H;
		io_rx_data = 512'hbfea23fffcafe3cf26e0eff20db3bacaccf8ebcb2a8e92f0fea2b00200b028be000000003fc823a3000000003453e9ee0000000031a5a1bd0000000048599232;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h31f0c0b810300e0cc33a9e3af3303eef723ba00c0c0038f930f38020030233f0000000003fc80a76000000003453c5a60000000031a59b8900000000485970db;#`PER_H;
		io_rx_data = 512'hbfea23fffcafe3cf26e0eff20db3bacaccf8ebcb2a8e92f0fea2b00200b028be000000003fc823a3000000003453e9ee0000000031a5a1bd0000000048599232;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hf2c3cfb8fe0cc87b0ef8dcfbcc3ca0f2ccbf08267cc3b0923ccf2f02f0aa0b3f000000003fc7e14c0000000034539fbb0000000031a598040000000048594d75;#`PER_H;
		io_rx_data = 512'h0030fc3300000c000080000000000000ab930000a0bdbf00c0af308070be000b000000003fc832ad000000003453f7e80000000031a5a358000000004859a793;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfef3ecccaff3cc32003cc8bbff3f3feacfbcb62ffaffe7bbe3c7fac3ba4bebac000000003fc75b3600000000345340c60000000031a58032000000004858dad2;#`PER_H;
		io_rx_data = 512'h0be3080b03df0fc3ef3d8bc2eb838be188efa80ce882702ca8ce6b8ecaabccbf000000003fc870e300000000345424550000000031a5af90000000004859de38;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hdfbffffecbff738bb3c9838bc20bc820ccbefc22fb9f0fc8fcc8cffc0efbfeff000000003fc4fde2000000003451a6740000000031a4fc39000000004856ddf1;#`PER_H;
		io_rx_data = 512'haaec30b0fff7aaaafb837f8cea2baa3c2f23fb3effefe00dfaf23af73328fb02000000003fc9d85f000000003454f3620000000031a5e56300000000485afbdc;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hdfbffffecbff738bb3c9838bc20bc820ccbefc22fb9f0fc8fcc8cffc0efbfeff000000003fc4fde2000000003451a6740000000031a4fc39000000004856ddf1;#`PER_H;
		io_rx_data = 512'h3ffffb3d20ffcfcacccffffffc3afcfcff2f0cc7f3ff83fffc7df3edfd8ffcef000000003fe26777000000003468ff750000000031ac1b4500000000486e24cf;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hfb3900332f32a02f3a200a823b230ecfea64ccf8cfbf3ca36ffffccfef4f7bfc000000003f7919ec000000003420df920000000031947fb200000000481c4ed0;#`PER_H;
		io_rx_data = 512'h3ffffb3d20ffcfcacccffffffc3afcfcff2f0cc7f3ff83fffc7df3edfd8ffcef000000003fe26777000000003468ff750000000031ac1b4500000000486e24cf;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'hffaaba0108e5c272338f07e0e38c78404a60b089c22da304d32902fb3f3c93fe000000003dfdcdae00000000333e817400000000313c1ea40000000046fee8ba;#`PER_H;
		io_rx_data = 512'h3ffffb3d20ffcfcacccffffffc3afcfcff2f0cc7f3ff83fffc7df3edfd8ffcef000000003fe26777000000003468ff750000000031ac1b4500000000486e24cf;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'h90b9130e2a044c5bfbbbb2a20a30acfccf6f3bffec38a22fecba0383893fcbfa000000003ab5f8d20000000030958dbd000000003091e974000000004362567d;#`PER_H;
		io_rx_data = 512'h3202b32b08033f08cebe80b773803c3f8f7f36ee33bbb31ef90fcc8fc03ffefc0000000041736d3d000000003583de3e0000000031f437490000000049e3a33c;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_data = 512'he8eccedcbecc0fbbe9cc8af1f5809048dfd7bb5fdefe5df6f5c3bffe3ffffe69000000002e38563c00000000265dfe18000000002e1ed23000000000362ca1fc;#`PER_H;
		io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;
		io_rx_rd_valid = 0; #150;#`PER_H;io_rx_rd_valid = 1;





		
		io_rx_rd_valid = 0;#`PER_H;
		
		#500;
		
		
		$finish; 
	end
	
	afu_core uut(
	.CLK_400M(CLK_400M),
    .reset_n(reset_n),
    
	//---------------------------------------------------
    //.spl_enable(spl_enable),
	.core_start(core_start),
	//---------------------------------------------------
	
    .spl_reset(spl_reset),
    
    // TX_RD request, afu_core --> afu_io
    .spl_tx_rd_almostfull(spl_tx_rd_almostfull),
    .cor_tx_rd_valid(cor_tx_rd_valid),
    .cor_tx_rd_addr(cor_tx_rd_addr),
    .cor_tx_rd_len(cor_tx_rd_len),  //[licheng]useless.
    
    
    // TX_WR request, afu_core --> afu_io
    .spl_tx_wr_almostfull(spl_tx_wr_almostfull),    
    .cor_tx_wr_valid(cor_tx_wr_valid),
    .cor_tx_dsr_valid(cor_tx_dsr_valid),
    .cor_tx_fence_valid(cor_tx_fence_valid),
    .cor_tx_done_valid(cor_tx_done_valid),
    .cor_tx_wr_addr(cor_tx_wr_addr), 
    .cor_tx_wr_len(cor_tx_wr_len), 
    .cor_tx_data(cor_tx_data),
             
    // RX_RD response, afu_io --> afu_core
    .io_rx_rd_valid(io_rx_rd_valid),
    .io_rx_data(io_rx_data),    
                 
    // afu_csr --> afu_core, afu_id
    .csr_id_valid(csr_id_valid),
    .csr_id_done(csr_id_done),    
    .csr_id_addr(csr_id_addr),
        
     // afu_csr --> afu_core, afu_ctx   
    .csr_ctx_base_valid(csr_ctx_base_valid),
    .csr_ctx_base(csr_ctx_base),

	.dsm_base_addr(dsm_base_addr),	
	.io_src_ptr(io_src_ptr),
	.io_dst_ptr(io_dst_ptr)

);

endmodule

