
`define CL 512
`define MAX_READ 64
`define READ_NUM_WIDTH 6
