
`define PER_H 2.5
`define PER_HH 1.25

module sim_afu_core();

	reg                             CLK_400M;
    reg                             reset_n;
    
	//---------------------------------------------------
    //reg                             spl_enable;
	reg 							core_start;
	//---------------------------------------------------
	
    reg                             spl_reset;
    
    // TX_RD request; afu_core --> afu_io
    reg                             spl_tx_rd_almostfull;
    wire                              cor_tx_rd_valid;
    wire  [57:0]                      cor_tx_rd_addr;
    wire  [5:0]                       cor_tx_rd_len;  //[licheng]useless.
    
    
    // TX_WR request; afu_core --> afu_io
    reg                             spl_tx_wr_almostfull;    
    wire                              cor_tx_wr_valid;
    wire                              cor_tx_dsr_valid;
    wire                              cor_tx_fence_valid;
    wire                              cor_tx_done_valid;
    wire  [57:0]                      cor_tx_wr_addr; 
    wire  [5:0]                       cor_tx_wr_len; 
    wire  [511:0]                     cor_tx_data;
             
    // RX_RD response; afu_io --> afu_core
    reg                             io_rx_rd_valid;
    reg [511:0]                     io_rx_data;    
                 
    // afu_csr --> afu_core; afu_id
    reg                             csr_id_valid;
    wire                              csr_id_done;    
    reg [31:0]                      csr_id_addr;
        
     // afu_csr --> afu_core; afu_ctx   
    reg                             csr_ctx_base_valid;
    reg [57:0]                      csr_ctx_base;

	reg  [63:0]	dsm_base_addr;	
	reg  [63:0] 						io_src_ptr;
	reg  [63:0] 						io_dst_ptr;
	
	//==========================
	//for test
	wire [6:0] backward_i_q_test; 
	wire [6:0] backward_j_q_test;
	
	//==========================
	
	initial forever #`PER_HH CLK_400M=!CLK_400M;
	
	always@(posedge CLK_400M)begin
	   if(cor_tx_rd_valid) begin
			
			$display("%h",cor_tx_rd_addr);
	   end
	end
	
	always@(*) $display("i = %h, j = %h\t",backward_i_q_test, backward_j_q_test);
	
//	always@(*) begin
//	   if(io_rx_rd_valid)
//	       $display("%h", io_rx_data);
	
//	end
	
	initial begin
		CLK_400M = 1;
		reset_n = 0;
		
		//---------------------------------------------------
		//spl_enable = 0;
		core_start = 0;
		//---------------------------------------------------
		
		spl_reset = 0;
		
		spl_tx_rd_almostfull = 0;
		spl_tx_wr_almostfull = 0;    

				 
		// RX_RD response = 0; afu_io --> afu_core
		io_rx_rd_valid = 0;
		io_rx_data = 0;    
					 
		// afu_csr --> afu_core = 0; afu_id
		csr_id_valid = 0;
		csr_id_addr = 0;
			
		 // afu_csr --> afu_core = 0; afu_ctx   
		csr_ctx_base_valid = 0;
		csr_ctx_base = 0;

		dsm_base_addr = 0;	
		io_src_ptr = 0;
		io_dst_ptr = 0;
		
		
		#0.1;
			
		#`PER_H;
		#`PER_H;
		
		reset_n = 1;
		
		#`PER_H;
		#`PER_H;
		
		core_start = 1;
		
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		
		io_rx_rd_valid = 1;
		io_rx_data[480] = 1; 
		io_rx_data[457:448] = 1; //batch size = 1;
		
		#`PER_H;
		
		io_rx_rd_valid = 0;
		io_rx_data = 0;
		
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#`PER_H;
		#300;
		io_rx_rd_valid = 1;

		io_rx_data = 512'h00000203030303020000020002000300010303030301030303030100000200030200020200000003010000010301010302030203020300020302010301000303;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000001020203030300030002020302000001020301030000020203020303030303010301020100;#`PER_H;
		io_rx_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea00000000000000001000000000000000f;#`PER_H;
		io_rx_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000010000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;
		
		io_rx_rd_valid = 0;
		
		#300;
        $display("%d",cor_tx_rd_valid);
		io_rx_rd_valid = 1; io_rx_data = 512'hc810c0030e0a8ec60220434000ca20e204c83c988f01c00c003c80018a042c8000000000182fb5f0000000001608a04a000000001a8f72c7000000002332667f;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he8eccedcbecc0fbbe9cc8af1f5809048dfd7bb5fdefe5df6f5c3bffe3ffffe69000000002e38563c00000000265dfe18000000002e1ed23000000000362ca1fc;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h550eff5ff77db4376975d17bdfccea5988e3269e22c92f30b3f93ffcdda9fbee00000000078b380d00000000072d0e630000000006e96251000000000d90bdbf;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h901177e582878f471e46ce4702db8e5061df340f812e20f987fcdc70dc1f6e3f000000000bdbf515000000000ad8057a000000000c7c48e70000000012fc5e0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb4c90339b30bd04a3ddea338f352443222ffe057fbbee1b7fc23bdbca13ff8f800000000307c76c7000000002831a9e7000000002e6a9acd0000000038f61b85;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4a82642e81bfc0cc8cccc0cf2c893bf0cc8ffefce80ba2f33bc88d41efbf02bf0000000031ab99f600000000290eed60000000002ea51c27000000003a5a2a83;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h213088a8cf0b0372ec220223b66208ccfeeb83f0233eb33cf2ecf00f2c020ff6000000003b4dfef600000000310bc1780000000030a5614200000000441450d0;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hebfca23c701c0800c01be31ada28a08e3b882cc809ecbc3f32e1d033c00efde7000000003b903a1d00000000314cf6700000000030b4063300000000445f7f40;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h643581088e499ac8517fcd32e2b21d619854c2d2973347cc895a3629cfdb5609000000000e83461b000000000e297a3f0000000010661a960000000017017590;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4c538155144c17c4b59481410c81a4b174e67204c75ff54ed091af7a0dc77474000000000e90692c000000000e3b4e8e00000000107b409000000000171886b6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h49b13cf3f1ef32e03b8ce88bcc0cfb0a2c40102cb00affcfcf2eee03ebef2a820000000032c53ae10000000029e79cee000000002ed7f538000000003b8675f9;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he2c06fc12be82b28c228c2bf0bcf9c2fffb3a2fbafedbacc020bbac0e08ef82c0000000032cb4bf30000000029ec8a80000000002ed926a4000000003b8c19e9;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfd03a14510c522c5fb7fbc0b56f714d5ffeee0ddc7f848ff35aff3246458f9ca0000000058b43c4a0000000042e3e0df000000003f70c244000000005d85bc93;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h364bdfd1f29f337b9f47f004d70ab484fd1eb7611206de1ff7116c578ee6c7b80000000058b5a0bc0000000042e56129000000003f726ab3000000005d8740e8;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4df3fccac8c1b4f33bfe6fdd7ee0c1f7d4d4c14e7e73dc3f4fa507df3dd5f3b300000000646f5f360000000049e464ac000000004909001a000000006720d984;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h2f8fefd7bebf7675b6d2367efef0ed27fcff85f9ff4ffcfb89bd5f3ba7f25e7100000000646fde570000000049e49ba0000000004909605b00000000672127ae;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc3f308eb38fcf3afefb33eef2a07eb0bfaffe3a03c1cff3f00ebf33ffbfe3cf3000000004786771b00000000393d3fb700000000331687a3000000004eebee8b;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h340af3f0ffcfeff8f0fc87f0fecffffffff0fffc9ccfbcfcfffff6334ecfffff000000004786895900000000393d51450000000033168a11000000004eebff51;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6ffd71870c7a67d464181121a9f6900a336c126ea34126843d5d900fdb3f41c100000000107cd8680000000010d571cd00000000139cdb500000000019fcc8fb;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h7086cc2b160700d2c140ff214041015805a18154806a8900d0018170e7cce57300000000107cdb810000000010d575e100000000139cdf2d0000000019fcce71;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdfc7124c81c420faffeb858c195f30fb08e234020082c81e4242ec50cd73ab09000000004ddbc265000000003cf0ef450000000036b65bd70000000054c32bff;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h74044481cca4e8fbfde44c2e665600038fe34c3afd88dc7c0cff443bfa850034000000004ddbc37a000000003cf0eff00000000036b65c810000000054c32d15;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'haaad2c088ff7ae6aaaaaaaaaaaaaaaaaabaaaaaaffaaaaaabf6ff87e7e267fee00000000604ebacb000000004841481200000000469fd6280000000064754afb;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6b73a14f547bc5b51f8f9fc06e3f0cfd7adedc6ea1a2ef07e371833e047c37cc00000000604ebb19000000004841487c00000000469fd6440000000064754b27;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc2c5d010d041036cf00039eeb78f33d5ef0a4d1185cdc37c23df60b49c7c3eff00000000675c04bb000000004b242037000000004aa951040000000068eea60a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h1f00b0f835c3f6ddfdc12daae0d9022dcb3ff0f8cc082bdf62cce5e2cdf3b10f00000000675c04e5000000004b242047000000004aa9511e0000000068eea636;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h2416f8e433a68f064c0bef1a2f0717990020c842f3f7373cafd57dcf5ee9ac2f000000002d693de10000000025f7290c000000002da2f5460000000035a024cd;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h2416f8e433a68f064c0bef1a2f0717990020c842f3f7373cafd57dcf5ee9ac2f000000002d693de10000000025f7290c000000002da2f5460000000035a024cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'ha8261d6de69b690be51dff05adab76d01ddce157f179e65fdef3aed69c222edd0000000024d8c499000000001fcd981e00000000261ef353000000002ed7d4f6;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'ha8261d6de69b690be51dff05adab76d01ddce157f179e65fdef3aed69c222edd0000000024d8c499000000001fcd981e00000000261ef353000000002ed7d4f6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcfff339f18f4505790b14613177af671f52c7b2b7710fe53976bf78f3f4cbd0000000054568f6f0000000040436eb1000000003bd5112c000000005a3316b4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcfff339f18f4505790b14613177af671f52c7b2b7710fe53976bf78f3f4cbd0000000054568f6f0000000040436eb1000000003bd5112c000000005a3316b4;#`PER_H;
		io_rx_rd_valid = 0; #500;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3810e3fff8020338f0f6e000ca0ac8fe20cc0f3efffffff2efcffffffffaecbf0000000043d6b8220000000036df3b4e000000003256f528000000004be1fbe8;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfe03fafca02fc33ffcafffcfef21f0433b03f88f74bfb800c04f3830be2c38c60000000043d6b93c0000000036df3bc2000000003256f53d000000004be1fcc5;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffffffffffffffffdfffffecfcfffe8acffcedf3ce0fff9b0f023f8cef2f0b0000000043d6b7c70000000036df3b40000000003256f525000000004be1fbd4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf33eff0334a3a3bf8363c1ece2b202faa0ef0ccb880206aa3f833b0a3320c0880000000043d6bef80000000036df3ec0000000003256f5fe000000004be200ca;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h00430cfd3e00ff0cc0ff30028ffb2f3a1ee23cfa33fb0f382fdff28ffefc38f00000000043d6a9780000000036df314b000000003256f2be000000004be1efff;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf33eff0334a3a3bf8363c1ece2b202faa0ef0ccb880206aa3f833b0a3320c0880000000043d6bef80000000036df3ec0000000003256f5fe000000004be200ca;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc0c880064b20b0fcf08033f0002dce03f3c9f04fffeccfcccf3bc8e3c5b0b36b0000000043d6796e0000000036df17fa000000003256ec95000000004be1c083;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h33f82cfcdff1836f37e00fff0f0008813c0333afcf3af02c0a1040ff0382f0c50000000043d70f280000000036df5ed100000000325702cb000000004be2323c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc0c880064b20b0fcf08033f0002dce03f3c9f04fffeccfcccf3bc8e3c5b0b36b0000000043d6796e0000000036df17fa000000003256ec95000000004be1c083;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h23c0fbecfb80c0efd832f2073233de9afbff2fce1c4f3fcf3df2fbcfe0cebebf0000000043d91b3a0000000036e04cba0000000032575feb000000004be387a1;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc0c880064b20b0fcf08033f0002dce03f3c9f04fffeccfcccf3bc8e3c5b0b36b0000000043d6796e0000000036df17fa000000003256ec95000000004be1c083;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3242f3e43cb238b4ffeec7dc8a23ac6880ff32bbc938efffaf0f720ef2f33fe40000000043de05f40000000036e2b9f90000000032587d63000000004be6d530;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc43fbff237fdffdf7f4d35cff53f777cde4543fe8fdffcc27cecf783ec93c300000000043d19c1f0000000036dc4fc30000000032561c0d000000004bdd1391;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcfffff335fbfffffe7fffadc4fc3fc1f3755f9fff3f7effffbcfffff64d0e2300000000043f038e80000000036ec690900000000325b6f1e000000004bf438f1;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf3fbff33fbef7f3dbf7f3ff3cfffffff3ffffff7effff0ff3f03f7ff8bcff5cc00000000439c718c0000000036bc92f60000000032494c0c000000004bacb5f2;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcfffff335fbfffffe7fffadc4fc3fc1f3755f9fff3f7effffbcfffff64d0e2300000000043f038e80000000036ec690900000000325b6f1e000000004bf438f1;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdf7ffcf7fe3ffffdc3f8bfcb03fcfcffeeb3e4c0ecf82fff31f33cbfccfcffc300000000432e42ce0000000036710ee000000000323691b2000000004b49ffa0;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h90830f80e3c31313cf220c3ecf0bbce2cff3fe3349220f1ac33cdb3fd3cff18c00000000448fb12300000000374d74b7000000003280f97b000000004c6cbaab;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3202b32b08033f08cebe80b773803c3f8f7f36ee33bbb31ef90fcc8fc03ffefc0000000041736d3d000000003583de3e0000000031f437490000000049e3a33c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he8eccedcbecc0fbbe9cc8af1f5809048dfd7bb5fdefe5df6f5c3bffe3ffffe69000000002e38563c00000000265dfe18000000002e1ed23000000000362ca1fc;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'ha9ed5556571bb57d55fad51551e6419659565d9579567455cc4655799bae6e750000000048c7c9310000000039ed5d8c000000003340e8a7000000004fd3521c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdd7946df41154ccf6c1a3e08aaaaaab1925ddaaaaaaaaaaeaaaaaaaaaacaaaaa000000005d11c6a400000000466cb8b9000000004463b2200000000061bde803;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'haaa3d676328be96ef84e6d4c021774e8494ab079d3a76fcd37d8768dfecde0b6000000005d11c6c600000000466cb91a000000004463b2680000000061bde838;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h342eb6aac2390ce80ef2ff23900c1145ba0815a23341207cd9860a7dfffffde2000000005d11c68000000000466cb89a000000004463b20b0000000061bde7db;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h7d571d9bd8eaaadc41e6f3339ce74c5555347201250087bc40549d336142d0b9000000005d11c83d00000000466cba74000000004463b4060000000061bde9c9;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h105bfc2810c5bc7b0c0c00c0d81802031803c099fce3f33e6f3575c0c8130e45000000005d11c37400000000466cb560000000004463ae050000000061bde427;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h7d571d9bd8eaaadc41e6f3339ce74c5555347201250087bc40549d336142d0b9000000005d11c83d00000000466cba74000000004463b4060000000061bde9c9;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd5178861d770f95f4f4cb356415e08612ff000197e5857d24575b518db3d1149000000005d11b7e800000000466cabca0000000044639f4e0000000061bdd800;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'haa07c33d0f7fa22800baf700fa142c008028d965fd35ea5f6348ff3ed3906c43000000005d11dc6100000000466cc551000000004463cf4c0000000061bdff82;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd5178861d770f95f4f4cb356415e08612ff000197e5857d24575b518db3d1149000000005d11b7e800000000466cabca0000000044639f4e0000000061bdd800;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6d489c84ccf1bb45f4ed8fe319bcd573ecfd3c43079e4295ce0405c87e50cdb1000000005d124b2900000000466d4d380000000044646c3c0000000061be77e3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd5178861d770f95f4f4cb356415e08612ff000197e5857d24575b518db3d1149000000005d11b7e800000000466cabca0000000044639f4e0000000061bdd800;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf11776ad00ba003cbe45d6e2fd90cef595475d972366f15ff195fcad8f2295f3000000005d1369a000000000466e629900000000446606b40000000061bf9493;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4757451d555d47955555e1f775555553659754d5ed9ffdea36c6ffb9371f0c0e000000005d10522600000000466bc9be00000000446259af0000000061bc87ed;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb88c55561cf053596d4c750ffe9c0c1dfd15f05c57c1f6257f348478cfdf6b53000000005d17e31b000000004671f35200000000446af0240000000061c4d36f;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h94f655015595456595d52d499de5554d96989597155dfc95bc131cc3dd70dd05000000005d03626100000000465f9e06000000004453e0060000000061aef293;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb88c55561cf053596d4c750ffe9c0c1dfd15f05c57c1f6257f348478cfdf6b53000000005d17e31b000000004671f35200000000446af0240000000061c4d36f;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5a64d56e66959605555655655b69e564554956555966567845559c586cfdfcaf000000005ce4ded500000000464bb5f10000000044352eba000000006191e100;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5cf537f57bdf5557f434d8136c9fd2c4cf2db436ac0ff6ccced782072c970125000000005d4044ae000000004691aa5b00000000449d9b760000000061e98801;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h75c15f7ff70e93bd5d5faea74abfdfcd7d9b672a8bfecec852f20554737d450d000000005c659f1a00000000460309e60000000043be88420000000061159d3e;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h01d565d96bc4fb55bcdf26551f5f7d51f7bde5d714ba55ea6167526d9fd77d52000000005e69721f00000000477bf8560000000045a642810000000063057d8a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5154d515bbfe9d55ffff2ffbfee3fbd7f671c3ff330f37bd33fdcc5ef37eed800000000057800f990000000041e911a9000000003e49e152000000005c4eb4ec;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h01d565d96bc4fb55bcdf26551f5f7d51f7bde5d714ba55ea6167526d9fd77d52000000005e69721f00000000477bf8560000000045a642810000000063057d8a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		
		spl_tx_rd_almostfull = 1;
		#2000;
		spl_tx_rd_almostfull = 0;
		
		
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6fadff5452c00182feb0322a8ef0cc2ffffff553fffefd55ffffffffffffffff000000004618cc1400000000387d9f000000000032de2bf3000000004dd9ea79;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6fadff5452c00182feb0322a8ef0cc2ffffff553fffefd55ffffffffffffffff000000004618cc1400000000387d9f000000000032de2bf3000000004dd9ea79;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffcffc40afddfcfbfee0283c2fdfffcf5f30cffd7fddffd7ffffd5d77ffbf000000004618cbc100000000387d9ef70000000032de2be1000000004dd9ea67;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3cfdc3ff3d2883f40e4f83bf870000ef7b4fb038fdd7d555c3ef1cf3aaac48ce000000004618ccbb00000000387d9f330000000032de2c1a000000004dd9eaf8;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h308c1130322c77062ff30eef30f30fe3f2fce0bc0ff30cccced2afdcc3cff8fc000000004618ca2600000000387d9e870000000032de2b99000000004dd9e9ba;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3cfdc3ff3d2883f40e4f83bf870000ef7b4fb038fdd7d555c3ef1cf3aaac48ce000000004618ccbb00000000387d9f330000000032de2c1a000000004dd9eaf8;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc8e4a3fff13c0bc0cfbeefff2ca1bcb0bc003bc0c020ec3ff98eae3ff0fcf3c3000000004618c67900000000387d9d3a0000000032de2b1f000000004dd9e5ae;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf7cf30cfff3ffea72f3fffef1cf7bb0b3cb8f3c3e3fc3faaf7c7302ff3c9303f000000004618d16000000000387da1530000000032de2cd5000000004dd9ee78;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc8e4a3fff13c0bc0cfbeefff2ca1bcb0bc003bc0c020ec3ff98eae3ff0fcf3c3000000004618c67900000000387d9d3a0000000032de2b1f000000004dd9e5ae;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcffff8ff02c4ffffffcf03ffffffbffeebfffbfcff0febcfff03f03e0efcfe00000000461919d500000000387db6cf0000000032de3836000000004dda0d26;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc8e4a3fff13c0bc0cfbeefff2ca1bcb0bc003bc0c020ec3ff98eae3ff0fcf3c3000000004618c67900000000387d9d3a0000000032de2b1f000000004dd9e5ae;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc30fc320bff23fbbdcfaf303ffbffbfccebbffcf2be9bf7be5fb83fffb33cac0000000004619a24d00000000387ded9a0000000032de4ba5000000004dda4f74;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0fc3383fce3d29f323c3fcbcfffef803fcb019cf333f03cce30f8402b7fcffe2000000004618667000000000387d71b60000000032de1a87000000004dd99fd3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf38c4083ef30d0b32f8f3ed0f13eff515ffd3dffcf8bf7ff3cabd3f8b0bcf69700000000461b250500000000387eb9a50000000032de905c000000004ddb4cfa;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5fffdffffffffef97ffffffd25efcfffc0bc5ccbf7ae0380868bfebb282c2f3b000000004612c04a00000000387b08ad0000000032dd029b000000004dd69aee;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf38c4083ef30d0b32f8f3ed0f13eff515ffd3dffcf8bf7ff3cabd3f8b0bcf69700000000461b250500000000387eb9a50000000032de905c000000004ddb4cfa;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcfffd57c57ffdd7f71f773dfddffff86cffdc701fffc7f3febbda3f2fb3cff00000000460aeecf00000000387633890000000032db9f8a000000004dd0bc9e;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffd4cf3f7f0decd31a8c8bf3ccddb1cf3cef0f43efeffc0de084dabf3ceafc000000004629505e000000003884eeb50000000032e1174c000000004de41ca1;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h7f74fe2383e3f6f3dcffafff3ef870bff2b1f20affc7e09b9a0b8afb0bcfffaf0000000045ea40f1000000003868053b0000000032d6a153000000004dbbeb01;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h83b3cf8cfbf07f3a34f3c6ff9cbcbfdf373ffc03a0bfcfb3fba0bf1bb63caaec0000000046966c170000000038b79d840000000032f0d815000000004e1edf50;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h90830f80e3c31313cf220c3ecf0bbce2cff3fe3349220f1ac33cdb3fd3cff18c00000000448fb12300000000374d74b7000000003280f97b000000004c6cbaab;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h83b3cf8cfbf07f3a34f3c6ff9cbcbfdf373ffc03a0bfcfb3fba0bf1bb63caaec0000000046966c170000000038b79d840000000032f0d815000000004e1edf50;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd0ba5147aa8455216d712557aab8aaaaaaaaaaaaaaaaaaaa5aaaaaa2a50ca925000000005d9d0dd50000000046e9c12700000000450a627a000000006250fc0a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd5557616d0256407aabb405675c2f60a4bb779c35de05d587425f555553db575000000005d9d0ddd0000000046e9c17300000000450a6296000000006250fc1a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd454957eff8ed155ce435038919d9b67009c6c2f54917d5d554b6545157d9445000000005d9d0d800000000046e9c09b00000000450a61bb000000006250fbaa;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd5557616d0256407aabb405675c2f60a4bb779c35de05d587425f555553db575000000005d9d0ddd0000000046e9c17300000000450a6296000000006250fc1a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h459bd9fd565ac057d5556185002f4e63eb9f7dcd53f45553c140d075d53d3ddd000000005d9d0ca10000000046e9c01c00000000450a6049000000006250fafa;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h10ecf1dc00d74d44b78ff456c45db5c7f4f56b319500614d7505646d1f554f35000000005d9d0ef00000000046e9c22000000000450a645e000000006250fd12;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h459bd9fd565ac057d5556185002f4e63eb9f7dcd53f45553c140d075d53d3ddd000000005d9d0ca10000000046e9c01c00000000450a6049000000006250fafa;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfc11ff7fb118f00c7b8400051141500d59414dc49f65fc5c355246073e34bdf1000000005d9d1ced0000000046e9c92700000000450a8f0600000000625105e6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h459bd9fd565ac057d5556185002f4e63eb9f7dcd53f45553c140d075d53d3ddd000000005d9d0ca10000000046e9c01c00000000450a6049000000006250fafa;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h58d5990af675d51db2f644f555bc9657455f13561eb18c3dd64c0933ddfcf45d000000005d9d57310000000046e9dab700000000450aba4100000000625117d7;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'had4d4fd6ef3477377c9ff7054045674cf730cdfbd54f58dd503355ff573af4bd000000005d9cf1a70000000046e9af4a00000000450a4094000000006250e67b;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h158083545415490b9e580739a1295de417d2d5dc5d5d5156dff06555ac5d4f62000000005d9db9f90000000046ea219100000000450b42810000000062516875;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h55d55554627e2b55977238b7ff4c37b34d36c3e3750ecc1f18bf3fc6177cff58000000005d9bd8000000000046e8caa5000000004507c9e900000000624fb4f2;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h158083545415490b9e580739a1295de417d2d5dc5d5d5156dff06555ac5d4f62000000005d9db9f90000000046ea219100000000450b42810000000062516875;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'haa855555e2c42b82afe6a99aef1922aeaba29eaaa6a2baead6eb89aa1bbbadca000000005d99ec610000000046e768670000000045057dac00000000624d7d8c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h8ef6721a004377c9835608cfe6d4d51c4c75cca4426977ab4afa4f4f22dca8ff000000005da148cf0000000046ed156e00000000450f4d7800000000625505cb;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf5d98577337d1535511543e3d9556547d5d71475565555d2461545d492afa786000000005d92389d0000000046ded0730000000044fe96d90000000062440297;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h510cd396bd2fd5555e708fc54905729fa4741525aaa5a682056beca53bfd6fe2000000005db66cd400000000471729a9000000004525df5d00000000626c57a6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5cf537f57bdf5557f434d8136c9fd2c4cf2db436ac0ff6ccced782072c970125000000005d4044ae000000004691aa5b00000000449d9b760000000061e98801;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h510cd396bd2fd5555e708fc54905729fa4741525aaa5a682056beca53bfd6fe2000000005db66cd400000000471729a9000000004525df5d00000000626c57a6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffaffbec8ce9b6eba95abc03555ffa77e69dc9beea8aaafff88a61d8d3c2300000000464bee2200000000389e15b10000000032e7698a000000004dfa1c23;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffaffbec8ce9b6eba95abc03555ffa77e69dc9beea8aaafff88a61d8d3c2300000000464bee2200000000389e15b10000000032e7698a000000004dfa1c23;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffaffbec8ce9b6eba95abc03555ffa77e69dc9beea8aaafff88a61d8d3c2300000000464bee2200000000389e15b10000000032e7698a000000004dfa1c23;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfff613f3e8d7a80f6fcc01ef09b88ef2f49aabe3fdfffcffffffffffffffffff00000000464bee5200000000389e15db0000000032e7699f000000004dfa1c34;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffaffbec8ce9b6eba95abc03555ffa77e69dc9beea8aaafff88a61d8d3c2300000000464bee2200000000389e15b10000000032e7698a000000004dfa1c23;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfff613f3e8d7a80f6fcc01ef09b88ef2f49aabe3fdfffcffffffffffffffffff00000000464bee5200000000389e15db0000000032e7699f000000004dfa1c34;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffaffbec8ce9b6eba95abc03555ffa77e69dc9beea8aaafff88a61d8d3c2300000000464bee2200000000389e15b10000000032e7698a000000004dfa1c23;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfff613f3e8d7a80f6fcc01ef09b88ef2f49aabe3fdfffcffffffffffffffffff00000000464bee5200000000389e15db0000000032e7699f000000004dfa1c34;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0ef8ea2f3c3fa0facc0e0d0f087be2eebb2cb4aa320f12f33eb82beeffcfe3ca00000000464bedf000000000389e158c0000000032e76986000000004dfa1bfe;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfff613f3e8d7a80f6fcc01ef09b88ef2f49aabe3fdfffcffffffffffffffffff00000000464bee5200000000389e15db0000000032e7699f000000004dfa1c34;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfe82cbff0030ff81a80bfc0bf0bc3befcf3fff7fcf60ff4dccbf37f83eeff08000000000464bedaf00000000389e15790000000032e76980000000004dfa1bd8;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heceffbb03fac2cf3cf3c0cd33f3b3f9fe810fb9ffce3f0038bb23182f8fe8ffc00000000464bee9f00000000389e15f00000000032e769a9000000004dfa1c48;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfe82cbff0030ff81a80bfc0bf0bc3befcf3fff7fcf60ff4dccbf37f83eeff08000000000464bedaf00000000389e15790000000032e76980000000004dfa1bd8;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hff000cf01fa0f0f03cf7fe2f533ff2b300eb3fd5f030c2bc23cd23330fef8cce00000000464bf1f600000000389e174f0000000032e76a3e000000004dfa1dfd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfe82cbff0030ff81a80bfc0bf0bc3befcf3fff7fcf60ff4dccbf37f83eeff08000000000464bedaf00000000389e15790000000032e76980000000004dfa1bd8;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcfb032ccbd3f3cfcfffe07c33e8fbdfcdf7ffbfdc71f00cffff3cbef0bfff2bc00000000464bfb0500000000389e1a680000000032e76b94000000004dfa21ff;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3e37ffcfc3c3ffa96873dac1afcef0ffffffaf1e033cb03cc3dfbeb73a7fdff100000000464be6ad00000000389e12a80000000032e768a7000000004dfa1604;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heef48354b0cc0340bfcc987ffebff63f6374f03fbdf2bff3cfc3ffe3f408303100000000464c1e3d00000000389e270d0000000032e77042000000004dfa3474;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h662b93faeff33fff3330373fcbffcfe403fb33030c3f2cfd833c3ef3fb262ea400000000464b7eba00000000389de3430000000032e74e34000000004df9e2cf;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heef48354b0cc0340bfcc987ffebff63f6374f03fbdf2bff3cfc3ffe3f408303100000000464c1e3d00000000389e270d0000000032e77042000000004dfa3474;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcffffffffbffdc33f7fcffeff3ffffcfbf0fffffffffffffefffffffffffffff00000000464ad58200000000389da5d40000000032e72f22000000004df98688;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hec3b0c0fc38ef3cffe7ef7f0fbfff3b3bcffd3f330fefc3f0eef30ffffceffff00000000464dcc1800000000389ea7770000000032e7a1b4000000004dfac8bd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heff3fe1e00084c2beff7ffb3ce3ce8c3feffeffdfbf3ffbffffffffffbffffff000000004645b46300000000389c5e350000000032e6b6a4000000004df7cfc4;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcfbfffffefffff3fffffbbffffffffffef7fffffffffbfbfffffffff7e3fff00000000466c325b0000000038a36e9c0000000032e98b3b000000004dffc5ce;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffffd4cf3f7f0decd31a8c8bf3ccddb1cf3cef0f43efeffc0de084dabf3ceafc000000004629505e000000003884eeb50000000032e1174c000000004de41ca1;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hffcfbfffffefffff3fffffbbffffffffffef7fffffffffbfbfffffffff7e3fff00000000466c325b0000000038a36e9c0000000032e98b3b000000004dffc5ce;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h9874a5d51751a52065869d3a18209194f5e17b3a58a01a9514b5609600000122000000005da7cbf00000000046f8a17d00000000451798c600000000625d49cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h9874a5d51751a52065869d3a18209194f5e17b3a58a01a9514b5609600000122000000005da7cbf00000000046f8a17d00000000451798c600000000625d49cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h9874a5d51751a52065869d3a18209194f5e17b3a58a01a9514b5609600000122000000005da7cbf00000000046f8a17d00000000451798c600000000625d49cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h0000000000000000000000000aaa9400902a8aa90a5dc15a580b872901adf343000000005da7cbe70000000046f8a16100000000451798b500000000625d4983;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h9874a5d51751a52065869d3a18209194f5e17b3a58a01a9514b5609600000122000000005da7cbf00000000046f8a17d00000000451798c600000000625d49cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4ac7cef43896c9975e223d76ba682306228c21572ee9ecbaaaaaad831eaaa8aa000000005da7cbce0000000046f8a12b000000004517989f00000000625d4968;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h9874a5d51751a52065869d3a18209194f5e17b3a58a01a9514b5609600000122000000005da7cbf00000000046f8a17d00000000451798c600000000625d49cd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4ac7cef43896c9975e223d76ba682306228c21572ee9ecbaaaaaad831eaaa8aa000000005da7cbce0000000046f8a12b000000004517989f00000000625d4968;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h957a62528a9965db2d2148aa7e7ffaa8ab6e5609778e52cb8a55541fee928368000000005da7cc6e0000000046f8a2510000000045179a4f00000000625d4a72;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4ac7cef43896c9975e223d76ba682306228c21572ee9ecbaaaaaad831eaaa8aa000000005da7cbce0000000046f8a12b000000004517989f00000000625d4968;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbe364c077dcdead59ab488fef3fe490aa8f15bcf8e3aaafeed34d75b5522bef7000000005da7ce660000000046f8a5120000000045179cff00000000625d4c09;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heaaa2e7bbe862a348fec8b27106913515f15b5f1a7e2ab85300248162dc586a6000000005da7ca640000000046f89f2b000000004517968e00000000625d47e3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heb8d25416c6a2f8fa98b7d909a6f1cd28d3059a2a9bd9f5a46a83ac7d1359aec000000005da7d5050000000046f8ae9a000000004517a8f100000000625d52f0;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6f26fc9317f64edcba5fe32c92a5f8e36bcafbccf1b033b2dfefc0d62ca5c809000000005da7b8470000000046f87e69000000004517753f00000000625d3411;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'heb8d25416c6a2f8fa98b7d909a6f1cd28d3059a2a9bd9f5a46a83ac7d1359aec000000005da7d5050000000046f8ae9a000000004517a8f100000000625d52f0;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h5555d58eaaaa99d5aeb2baaaaaaaaeaaaeaa8aaaaaaaaaaaaa8a2abaa68baaa8000000005da793490000000046f84f5e00000000451745af00000000625d0eaa;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb7366aad6e9ebeb926a5de9269d02ae4d87ab26feb1a5870bba4cea65addb1e2000000005da81d250000000046f9538d00000000451804d900000000625db7f5;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h8e534ba348c4a22a9d01234479cde4c8b12f12dcae1c3b95e6eaee3aabaefbe2000000005da6d90c0000000046f5d5e4000000004516a9f100000000625bbd1f;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h55d15355713d74d5eed50f5deeaaebe7acc6a6adae8ae66aabb9abfabab6ea62000000005daae2aa00000000470ecdc000000000451a7c5a000000006261673c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h8ef6721a004377c9835608cfe6d4d51c4c75cca4426977ab4afa4f4f22dca8ff000000005da148cf0000000046ed156e00000000450f4d7800000000625505cb;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h55d15355713d74d5eed50f5deeaaebe7acc6a6adae8ae66aabb9abfabab6ea62000000005daae2aa00000000470ecdc000000000451a7c5a000000006261673c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hec2900f2d61d3f1ff7f351dd09c377d4e5c3d755198fff441fbfdf73016c5c2700000000155a6ece00000000146be1990000000018443d6c000000002052bb2d;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'he5c3c7c7cf205997a2aa49e4aaa9aaaaaaaaaaaaaaaaa6aa8aaa62aad44cf52000000000155a6efe00000000146be1a50000000018443d91000000002052bb4c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hec2900f2d61d3f1ff7f351dd09c377d4e5c3d755198fff441fbfdf73016c5c2700000000155a6ece00000000146be1990000000018443d6c000000002052bb2d;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h4a518f14099c324bdd621c9906726d05b46925fe65db504b3d794ae5cb8ba2a800000000155a6f0e00000000146be1ee0000000018443da5000000002052bb5f;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hec2900f2d61d3f1ff7f351dd09c377d4e5c3d755198fff441fbfdf73016c5c2700000000155a6ece00000000146be1990000000018443d6c000000002052bb2d;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf4047445a33b9edf479c95151bd43109b21eabfd6a7bb926772be8dff700938b00000000155a6f7e00000000146be2660000000018443e39000000002052bbe3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h58f37b1d44c95557f7f52436fd5dffbdc7d753e37515fd5cd9954dd55555555d00000000155a6e3e00000000146be1670000000018443cf2000000002052bae9;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc0331f9dbb7f034f444cdf99cb051b180226417acf000105b318f70f0238d44200000000155a71f100000000146be37a0000000018444004000000002052bd91;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf3d781b2e9377809344b9cf5d05c234a830485c6c3f2815e0950008fa4ccdb8000000000155a699600000000146bdcdf0000000018443768000000002052b623;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hc0331f9dbb7f034f444cdf99cb051b180226417acf000105b318f70f0238d44200000000155a71f100000000146be37a0000000018444004000000002052bd91;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdd886457f0bf2ccb30eb7fc4bd001337404c8778df7fd31f1ffff3dc173ff3ff00000000155a5e3300000000146bd5160000000018442fe5000000002052ab52;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb19833347ef2403b042dd6c71e8423cc0f37d2b5bdef5df0775edd08d2d0793700000000155aacef00000000146bee4d0000000018445113000000002052cbb1;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbecbccfc0df90dcdf4f044ffcf067719bc13d7fd9b733933cd4e04b5ec53e35f000000001559ad1800000000146bb14c000000001843ebd900000000205272c3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3401fa052070043780a2874a0e0ecafb3314c7074bc6738fc37c24f12fcb37ec00000000155c71e600000000146c5b450000000018451ebb0000000020537b1a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h22e0c8d01d13e8161d07c1dc4d7ce67176b1514d3355150b41553cefe35fd076000000001557cb4d00000000146a2c49000000001842577b000000002050b66f;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3401fa052070043780a2874a0e0ecafb3314c7074bc6738fc37c24f12fcb37ec00000000155c71e600000000146c5b450000000018451ebb0000000020537b1a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc3ffbc8cbcbb827338e3afcc737efa00aa3e0fffff3ff0b555555df555555550000000034c73d21000000002ba894c6000000002f3b22c7000000003da2b5d2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc3ffbc8cbcbb827338e3afcc737efa00aa3e0fffff3ff0b555555df555555550000000034c73d21000000002ba894c6000000002f3b22c7000000003da2b5d2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc3ffbc8cbcbb827338e3afcc737efa00aa3e0fffff3ff0b555555df555555550000000034c73d21000000002ba894c6000000002f3b22c7000000003da2b5d2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc3ffbc8cbcbb827338e3afcc737efa00aa3e0fffff3ff0b555555df555555550000000034c73d21000000002ba894c6000000002f3b22c7000000003da2b5d2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc3ffbc8cbcbb827338e3afcc737efa00aa3e0fffff3ff0b555555df555555550000000034c73d21000000002ba894c6000000002f3b22c7000000003da2b5d2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h03e8f3003c2832ce83faffa02a02e3ce88f38fcc8c3c0ebcc2af887eaeaaaaa80000000034c73d53000000002ba894da000000002f3b22e7000000003da2b5ec;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd57fff5de33e3ea23fe83f03233c7afa9f5bf00d20287eafed220ebc82fc23c80000000034c73cf0000000002ba894a8000000002f3b22b9000000003da2b5af;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'habaaaaaa383eaaaa238fca2b08b80ceec3fc39c8ca0f803cbfe83c2bc300b0f80000000034c73d9d000000002ba89533000000002f3b22ed000000003da2b643;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h00c0200ba3a1f32030a82ea0cc3b00ba0bebc8bcfee123d03b08382ef3cbc01c0000000034c73be8000000002ba8927e000000002f3b2297000000003da2b483;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'habaaaaaa383eaaaa238fca2b08b80ceec3fc39c8ca0f803cbfe83c2bc300b0f80000000034c73d9d000000002ba89533000000002f3b22ed000000003da2b643;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h2f08c0fe0200f3b3fcaf33ebf81bf28ab33fc8fc23888f28e23f8808000c0fc00000000034c739a0000000002ba89109000000002f3b20a1000000003da2b236;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3028aacca0093ea02f3013f08f73fbbc2d33fbe83323c0f2ceb4eb0f3a03f0c30000000034c74110000000002ba89952000000002f3b235c000000003da2b942;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h30fbfafee3cf723ccfea48ff800a8d8a2308308cb03c2f3ec832032f38cb207c0000000034c72bd1000000002ba88870000000002f3b1fc8000000003da2a5f7;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h82ffe81cf3f37c83c028cfbe0f2f2e3bacd8dfc3e8a4f00db8c3f0c8c30f000e0000000034c76635000000002ba8b80c000000002f3b2894000000003da2dd2b;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3f8c283202fbc20b033220c3f3f680fcc88cbff337028f3f7fcec20f8fffc1bf0000000034c695ac000000002ba83886000000002f3b0f35000000003da21799;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h82ffe81cf3f37c83c028cfbe0f2f2e3bacd8dfc3e8a4f00db8c3f0c8c30f000e0000000034c76635000000002ba8b80c000000002f3b2894000000003da2dd2b;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3572f4a103e3a5ef52fad371b512f6e1696ef7e5aaaaaaaa2d6f57ba465fcb5c000000005931b9ab0000000043550ca9000000003fffbb79000000005e0a1cb3;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb80dee6413d6603cea927e26a47345588ba44297bfc4fec21066f064d799669d000000005931b9cd0000000043550cd3000000003fffbb9b000000005e0a1cc5;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbaae08a2ef28a2226873acbcddad0d6d3d2aa0624b6932b8a78c8fcd39022c2e000000005931b9430000000043550c43000000003fffbb22000000005e0a1c58;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hb80dee6413d6603cea927e26a47345588ba44297bfc4fec21066f064d799669d000000005931b9cd0000000043550cd3000000003fffbb9b000000005e0a1cc5;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h960ce3305c218e3efff89e882fc12a0b608ec19ee8eaee00818fa9d9bfff69a4000000005931b8dc0000000043550b81000000003fffbac3000000005e0a1be0;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h6dfc04c582ffd5db41a30554da0caf6888c250e60ac11939cfa09f1bfbfabc2b000000005931ba910000000043550df2000000003fffbc57000000005e0a1da6;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'ha8e796027a063383de039afeabac6713fe8961e1673286aabeaea9d8abaffaf4000000005931b6340000000043550511000000003fffb8d5000000005e0a18e6;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd699b2cd91e4d0c4dbdcc3e755f949d83a215ba57f8fb5ffbd4129b168eaaf1b000000005931c23b0000000043551a28000000003fffc554000000005e0a25c9;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfd0f483d30dde71e6607d43001b98f187acca28e88bbd2096a6d05d6f319ef000000000059319dab000000004354ba1e000000003fff9e87000000005e0a00b0;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd699b2cd91e4d0c4dbdcc3e755f949d83a215ba57f8fb5ffbd4129b168eaaf1b000000005931c23b0000000043551a28000000003fffc554000000005e0a25c9;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbfffffff810cccf3eea083bfaaeee00f30efafa28c40000c37f3f0e03eb0b0c8000000004506d9990000000037a8188500000000329e583d000000004ce98aa5;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf020030bfe62e100feb2fbb0cacf233b2ffea26dc70e81e0cec08ce6ff5cf27f000000004506d9ce0000000037a818a000000000329e5840000000004ce98ad2;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h18200b7dea82e10bfcff1f3cffcb1febffffff1f3fffffffff0efc8effffffff000000004506d92b0000000037a8185f00000000329e5832000000004ce98a44;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hea7fc1cdbf3f8b8fbfff224330f0cdb3f043203820f83dffffcccff8fffabcff000000004506da300000000037a818f100000000329e584c000000004ce98b13;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hbf3fcfd0fef3ffbc8eff370ff30efaaffaffffffffffffffef35dff32ca4abeb000000004506d4510000000037a817c800000000329e5808000000004ce9895f;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf21dfcf88022fab00f0eabb32cfbcceffffc04ffffff75ffeffcff3fbf00b2ff000000004506e1d80000000037a81ac100000000329e58ad000000004ce98d3a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hcc33ff0ba1f3f30c30f90000f08330bfffcbf8e0dfaa033f3ecfb3f2fa33fff80000000045069c830000000037a80e0300000000329e56a0000000004ce9815a;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf21dfcf88022fab00f0eabb32cfbcceffffc04ffffff75ffeffcff3fbf00b2ff000000004506e1d80000000037a81ac100000000329e58ad000000004ce98d3a;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h3d9ac618ca900f0a8003cf2f0081d14ccd49180fae1fffff3fc78916ab382c850000000026144973000000002100e652000000002776212f00000000300d370c;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h082bbfffc05022dbb0c84f89cf7c7badb7117606f53453f1fbad62182b5ec0420000000026144998000000002100e66d000000002776214300000000300d3738;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h82ffa76b2383b10d5e2908899032ad5946f201853aad6c3b382e05332680180200000000261448bd000000002100e61100000000277620f700000000300d36bb;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h082bbfffc05022dbb0c84f89cf7c7badb7117606f53453f1fbad62182b5ec0420000000026144998000000002100e66d000000002776214300000000300d3738;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hf1bdc2dd3fffffff5fffcd6f8083fcfcffff7fb1fffffffff9ffffffffffffff0000000054ac18fa00000000407dd83e000000003c38b36e000000005a7b05da;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfffffffffffffcff1fe7beff01cf8f403f9d804ac3fa36bdfe53528de00fd3e70000000054ac18b500000000407dd82d000000003c38b35e000000005a7b05c0;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'h51cdc4df04b605ee5555555bd55555552560393047fe2fcef75b54d5f2fffffe0000000054ac195b00000000407dd845000000003c38b379000000005a7b05e7;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd6c49b47737554512e56147a0506bcc1d2559f77601f1d6b555169695575946900000000290190650000000022ecb3590000000029ed4b07000000003257543b;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd6c49b47737554512e56147a0506bcc1d2559f77601f1d6b555169695575946900000000290190650000000022ecb3590000000029ed4b07000000003257543b;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd6c49b47737554512e56147a0506bcc1d2559f77601f1d6b555169695575946900000000290190650000000022ecb3590000000029ed4b07000000003257543b;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdfb3720e50cd4324b349ffd2ff0e50081f6dffff57f851ba5555555555455555000000002901907b0000000022ecb36f0000000029ed4b440000000032575452;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hd6c49b47737554512e56147a0506bcc1d2559f77601f1d6b555169695575946900000000290190650000000022ecb3590000000029ed4b07000000003257543b;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hdfb3720e50cd4324b349ffd2ff0e50081f6dffff57f851ba5555555555455555000000002901907b0000000022ecb36f0000000029ed4b440000000032575452;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 0; #200;;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 1; io_rx_data = 512'hfed905783dc5548e2257bbf361041750105690d05de78f1236014003a1409d54000000000af9cfdd000000000a1c9378000000000b50e7ae0000000011f008fd;#`PER_H;
		io_rx_rd_valid = 0; #200;

		
		#5000;
		
		
		$finish; 
	end
	
	afu_core uut(
	.CLK_400M(CLK_400M),
    .reset_n(reset_n),
    
	//---------------------------------------------------
    //.spl_enable(spl_enable),
	.core_start(core_start),
	//---------------------------------------------------
	
    .spl_reset(spl_reset),
    
    // TX_RD request, afu_core --> afu_io
    .spl_tx_rd_almostfull(spl_tx_rd_almostfull),
    .cor_tx_rd_valid(cor_tx_rd_valid),
    .cor_tx_rd_addr(cor_tx_rd_addr),
    .cor_tx_rd_len(cor_tx_rd_len),  //[licheng]useless.
    
    
    // TX_WR request, afu_core --> afu_io
    .spl_tx_wr_almostfull(spl_tx_wr_almostfull),    
    .cor_tx_wr_valid(cor_tx_wr_valid),
    .cor_tx_dsr_valid(cor_tx_dsr_valid),
    .cor_tx_fence_valid(cor_tx_fence_valid),
    .cor_tx_done_valid(cor_tx_done_valid),
    .cor_tx_wr_addr(cor_tx_wr_addr), 
    .cor_tx_wr_len(cor_tx_wr_len), 
    .cor_tx_data(cor_tx_data),
             
    // RX_RD response, afu_io --> afu_core
    .io_rx_rd_valid(io_rx_rd_valid),
    .io_rx_data(io_rx_data),    
                 
    // afu_csr --> afu_core, afu_id
    .csr_id_valid(csr_id_valid),
    .csr_id_done(csr_id_done),    
    .csr_id_addr(csr_id_addr),
        
     // afu_csr --> afu_core, afu_ctx   
    .csr_ctx_base_valid(csr_ctx_base_valid),
    .csr_ctx_base(csr_ctx_base),

	.dsm_base_addr(dsm_base_addr),	
	.io_src_ptr(io_src_ptr),
	.io_dst_ptr(io_dst_ptr),
	
	.backward_i_q_test(backward_i_q_test), 
	.backward_j_q_test(backward_j_q_test)

);

endmodule

